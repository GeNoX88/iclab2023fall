//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Fall
//   Lab01 Exercise		: Supper MOSFET Calculator
//   Author     		: Lin-Hung Lai (lhlai@ieee.org)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : SMC.v
//   Module Name : SMC
//   Release version : V1.0 (Release Date: 2023-09)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

// my best is 38732
module SMC (
  input [2:0] W_0,  //    1~7 unsigned integer
  input [2:0] V_GS_0,  // 1~7 unsigned integer
  input [2:0] V_DS_0,  // 1~7 unsigned integer
  input [2:0] W_1,  //    1~7 unsigned integer
  input [2:0] V_GS_1,  // 1~7 unsigned integer
  input [2:0] V_DS_1,  // 1~7 unsigned integer
  input [2:0] W_2,  //    1~7 unsigned integer
  input [2:0] V_GS_2,  // 1~7 unsigned integer
  input [2:0] V_DS_2,  // 1~7 unsigned integer
  input [2:0] W_3,  //    1~7 unsigned integer
  input [2:0] V_GS_3,  // 1~7 unsigned integer
  input [2:0] V_DS_3,  // 1~7 unsigned integer
  input [2:0] W_4,  //    1~7 unsigned integer
  input [2:0] V_GS_4,  // 1~7 unsigned integer
  input [2:0] V_DS_4,  // 1~7 unsigned integer
  input [2:0] W_5,  //    1~7 unsigned integer
  input [2:0] V_GS_5,  // 1~7 unsigned integer
  input [2:0] V_DS_5,  // 1~7 unsigned integer
  input [1:0] mode, //    mode[1]==1'b1...larger, mode[1]==1'b0...smaller; mode[0]==1'b1...weighted avg I(*3,*4,*5,/12); mode[0]==1'b0...avg g(*1,*1,*1,/3)
  output [7:0] out_n  // 0~255 unsigned integer (an avg number)
);
  integer i, j;
  wire [2:0] W[0:5];
  wire [2:0] V_GS[0:5];
  wire [2:0] V_DS[0:5];
  assign W[0] = W_0;
  assign W[1] = W_1;
  assign W[2] = W_2;
  assign W[3] = W_3;
  assign W[4] = W_4;
  assign W[5] = W_5;

  assign V_GS[0] = V_GS_0;
  assign V_GS[1] = V_GS_1;
  assign V_GS[2] = V_GS_2;
  assign V_GS[3] = V_GS_3;
  assign V_GS[4] = V_GS_4;
  assign V_GS[5] = V_GS_5;

  assign V_DS[0] = V_DS_0;
  assign V_DS[1] = V_DS_1;
  assign V_DS[2] = V_DS_2;
  assign V_DS[3] = V_DS_3;
  assign V_DS[4] = V_DS_4;
  assign V_DS[5] = V_DS_5;


  reg [2:0] V_on[0:5];
  reg region[0:5];

  always @(*) begin
    for (i = 0; i < 6; i = i + 1) begin
      V_on[i]   = V_GS[i] - 1;  // V_on = 0~6
      region[i] = V_on[i] > V_DS[i];
    end
  end

  // region:
  //  if(V_on > V_DS) -> (6, 5)~(6,1), (5,4)~(5,1), (4,3)~(4,1), (3,2)~(3,1), (2,1)
  //    I = (1/3)[W(2*V_on*V_DS-V_DS^2)] = [W*V_DS(2*V_on-V_DS)]/3
  //      min = 3/3 = 1
  //      max at V_on=6, V_DS=5, max = (1/3)*7*5*7 = 245/3 8bit=>7bit
  //    g = (W*V_DS*2)/3
  //      min = 2/3 = 0
  //      max = (2/3)*7*7 = 98/3 7bit=>6bit
  //  if(V_on <= V_DS) -> (66~67), (55~57), (44~47), (33~37), (22~27), (11~17), (01~07)
  //    I = (W*V_on^2)/3
  //      min = 0
  //      max = (1/3)*7*36 = 252/3=84 8bit=>7bit
  //    g = (W*V_on * 2)/3
  //      min = 0
  //      max = (2/3)*7*6 = 84/3=26 7bit=>6bit

  //************ 8 bit prototype ************************
  reg [7:0] Ig[0:5];
  wire [7:0] a[0:5];
  wire [7:0] b[0:5];
  wire [7:0] c[0:5];
  wire [7:0] d[0:5];
  wire [7:0] e[0:5];


  //******* cell area smallest *******************
  reg [2:0] V[0:5];
  reg [4:0] B[0:5];
  always @(*) begin
    for (j = 0; j < 6; j = j + 1) begin
      V[j]  = region[j] ? V_DS[j] : V_on[j];
      B[j]  = ~mode[0] ? 2 : region[j] ? ((V_on[j] << 1) - V_DS[j]) : V_on[j];
      Ig[j] = W[j] * V[j] * B[j];
    end
  end
  //*************************************************

  wire cmp[0:11];
  assign cmp[0] = Ig[0] > Ig[4];
  assign cmp[1] = Ig[1] > Ig[5];
  assign cmp[2] = Ig[2] > Ig[3];
  assign cmp[3] = a[0] > a[5];
  assign cmp[4] = a[1] > a[2];
  assign cmp[5] = a[3] > a[4];
  assign cmp[6] = b[0] > b[1];
  assign cmp[7] = b[2] > b[3];
  assign cmp[8] = b[4] > b[5];
  assign cmp[9] = c[1] > c[2];
  assign cmp[10] = c[3] > c[4];
  assign cmp[11] = d[2] > d[3];

  // the "smallest" one of optimal sorting networks
  // [[1 5][2 6][3 4][1 6][2 3][4 5][1 2][3 4][5 6][2 3][4 5][3 4]]
  assign {a[0], a[4]} = cmp[0] ? {Ig[0], Ig[4]} : {Ig[4], Ig[0]};
  assign {a[1], a[5]} = cmp[1] ? {Ig[1], Ig[5]} : {Ig[5], Ig[1]};
  assign {a[2], a[3]} = cmp[2] ? {Ig[2], Ig[3]} : {Ig[3], Ig[2]};
  assign {b[0], b[5]} = cmp[3] ? {a[0], a[5]} : {a[5], a[0]};
  assign {b[1], b[2]} = cmp[4] ? {a[1], a[2]} : {a[2], a[1]};
  assign {b[3], b[4]} = cmp[5] ? {a[3], a[4]} : {a[4], a[3]};
  assign {c[0], c[1]} = cmp[6] ? {b[0], b[1]} : {b[1], b[0]};
  assign {c[2], c[3]} = cmp[7] ? {b[2], b[3]} : {b[3], b[2]};
  assign {c[4], c[5]} = cmp[8] ? {b[4], b[5]} : {b[5], b[4]};
  assign {d[1], d[2]} = cmp[9] ? {c[1], c[2]} : {c[2], c[1]};
  assign {d[3], d[4]} = cmp[10] ? {c[3], c[4]} : {c[4], c[3]};
  assign {e[2], e[3]} = cmp[11] ? {d[2], d[3]} : {d[3], d[2]};


  wire [7:0] n0 = c[0], n1 = d[1], n2 = e[2], n3 = e[3], n4 = d[4], n5 = c[5];


  wire [7:0] MOS1_3x, MOS2_3x, MOS3_3x;  // 0~252 8bit 
  wire [6:0] MOS1, MOS2, MOS3;  // 0~84 7bit
  assign {MOS1_3x, MOS2_3x, MOS3_3x} = mode[1] ? {n0, n1, n2} : {n3, n4, n5};

  divider_3_LUT MOS1_ (
    MOS1_3x,
    MOS1
  );
  divider_3_LUT MOS2_ (
    MOS2_3x,
    MOS2
  );
  divider_3_LUT MOS3_ (
    MOS3_3x,
    MOS3
  );
  // // ************* prototype *******************
  // assign out_n = mode[0] ?
  //     // (MOS1 * 3 + MOS2 * 4 + MOS3 * 5) / 12 :
  //     // (MOS1 * 3 + MOS3 * 5 + MOS2 * 4) / 12:
  //     // (MOS2 * 4+MOS1 * 3 + MOS3 * 5  ) / 12:
  //     (MOS2 * 4 + MOS3 * 5 + MOS1 * 3) / 12 :  // V
  //     // (MOS3 * 5+MOS1 * 3 +  + MOS2 * 4) / 12:
  //     // (MOS3 * 5+MOS2 * 4+MOS1 * 3  ) / 12:
  //     // (MOS1 + MOS2 + MOS3) / 3;  // 26235 combinations
  //     // (MOS1 + MOS3 + MOS2) / 3;  // 26235 combinations
  //     (MOS2 + MOS1 + MOS3) / 3;  // 26235 combinations V
  // // (MOS2 + MOS3 + MOS1) / 3;  // 26235 combinations
  // // (MOS3 + MOS1 + MOS2) / 3;  // 26235 combinations
  // // (MOS3 + MOS2 + MOS1) / 3;  // 26235 combinations
  // // **************************************************

  // ******** Lin's solution(smallest area solution - 38732) *****************

  wire [9:0] total_4x = mode[0]?
    ((MOS2<<2)+((MOS3<<2)+MOS3)+((MOS1<<1)+MOS1)) :
      ((MOS2<<2)+(MOS1<<2)+((MOS3<<2)));

  wire [6:0] out_7bit;
  divider_12_LUT TOTAL (
    total_4x,
    out_7bit
  );
  assign out_n = {1'b0, out_7bit};

  // ********** replace //12 with //4 then //3 ****************************
  // wire [6:0] out_7bit;
  // assign out_n = {1'b0, out_7bit};
  // wire [7:0] out_3x = mode[0]? 
  // ((MOS3 * 5 + MOS1 * 3)/4 + MOS2):
  // (MOS2 + MOS1 + MOS3);
  // divider_3_LUT OUT_N (
  //   out_3x,
  //   out_7bit
  // );

  // ******************************************
endmodule



module divider_12_ning (
  input [9:0] dividend,  // 0~1023
  output reg [6:0] q
);
  always @(*) begin
    q = (dividend*((1<<9)+(1<<7)+(1<<5)+(1<<3)+(1<<1)+1)) >> 13;
  end
endmodule
module divider_3_ning (
  input [7:0] dividend,  // 0~252
  output reg [6:0] q
);
  wire [14:0] high = 
  (dividend << 7) + (dividend << 5) + (dividend << 3 ) + (dividend << 1) + (dividend << 0);
  always @(*) begin
    q = high >> 9;
  end
endmodule

module divider_3_LUT (
  input [7:0] dividend,  // 0~255
  output reg [6:0] q  // 0~84 7bit
);
  always @(*) begin
    case (dividend)
      0, 1, 2: q = 0;
      3, 4, 5: q = 1;
      6, 7, 8: q = 2;
      9, 10, 11: q = 3;
      12, 13, 14: q = 4;
      15, 16, 17: q = 5;
      18, 19, 20: q = 6;
      21, 22, 23: q = 7;
      24, 25, 26: q = 8;
      27, 28, 29: q = 9;
      30, 31, 32: q = 10;
      33, 34, 35: q = 11;
      36, 37, 38: q = 12;
      39, 40, 41: q = 13;
      42, 43, 44: q = 14;
      45, 46, 47: q = 15;
      48, 49, 50: q = 16;
      51, 52, 53: q = 17;
      54, 55, 56: q = 18;
      57, 58, 59: q = 19;
      60, 61, 62: q = 20;
      63, 64, 65: q = 21;
      66, 67, 68: q = 22;
      69, 70, 71: q = 23;
      72, 73, 74: q = 24;
      75, 76, 77: q = 25;
      78, 79, 80: q = 26;
      81, 82, 83: q = 27;
      84, 85, 86: q = 28;
      87, 88, 89: q = 29;
      90, 91, 92: q = 30;
      93, 94, 95: q = 31;
      96, 97, 98: q = 32;
      99, 100, 101: q = 33;
      102, 103, 104: q = 34;
      105, 106, 107: q = 35;
      108, 109, 110: q = 36;
      111, 112, 113: q = 37;
      114, 115, 116: q = 38;
      117, 118, 119: q = 39;
      120, 121, 122: q = 40;
      123, 124, 125: q = 41;
      126, 127, 128: q = 42;
      129, 130, 131: q = 43;
      132, 133, 134: q = 44;
      135, 136, 137: q = 45;
      138, 139, 140: q = 46;
      141, 142, 143: q = 47;
      144, 145, 146: q = 48;
      147, 148, 149: q = 49;
      150, 151, 152: q = 50;
      153, 154, 155: q = 51;
      156, 157, 158: q = 52;
      159, 160, 161: q = 53;
      162, 163, 164: q = 54;
      165, 166, 167: q = 55;
      168, 169, 170: q = 56;
      171, 172, 173: q = 57;
      174, 175, 176: q = 58;
      177, 178, 179: q = 59;
      180, 181, 182: q = 60;
      183, 184, 185: q = 61;
      186, 187, 188: q = 62;
      189, 190, 191: q = 63;
      192, 193, 194: q = 64;
      195, 196, 197: q = 65;
      198, 199, 200: q = 66;
      201, 202, 203: q = 67;
      204, 205, 206: q = 68;
      207, 208, 209: q = 69;
      210, 211, 212: q = 70;
      213, 214, 215: q = 71;
      216, 217, 218: q = 72;
      219, 220, 221: q = 73;
      222, 223, 224: q = 74;
      225, 226, 227: q = 75;
      228, 229, 230: q = 76;
      231, 232, 233: q = 77;
      234, 235, 236: q = 78;
      237, 238, 239: q = 79;
      240, 241, 242: q = 80;
      243, 244, 245: q = 81;
      246, 247, 248: q = 82;
      249, 250, 251: q = 83;
      252, 253, 254: q = 84;
      255: q = 85;
      default: q = 8'dx;
    endcase
  end
endmodule
module divider_12_LUT (
  input [9:0] dividend,  // 0~1023
  output reg [6:0] q
);
  always @(*) begin
    case (dividend)
      0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11: q = 0;
      12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23: q = 1;
      24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35: q = 2;
      36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47: q = 3;
      48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59: q = 4;
      60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71: q = 5;
      72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83: q = 6;
      84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95: q = 7;
      96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 107: q = 8;
      108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119: q = 9;
      120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131: q = 10;
      132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143: q = 11;
      144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155: q = 12;
      156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167: q = 13;
      168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179: q = 14;
      180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191: q = 15;
      192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203: q = 16;
      204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215: q = 17;
      216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227: q = 18;
      228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239: q = 19;
      240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251: q = 20;
      252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263: q = 21;
      264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275: q = 22;
      276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287: q = 23;
      288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299: q = 24;
      300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311: q = 25;
      312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323: q = 26;
      324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335: q = 27;
      336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347: q = 28;
      348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359: q = 29;
      360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371: q = 30;
      372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383: q = 31;
      384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395: q = 32;
      396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 407: q = 33;
      408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419: q = 34;
      420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431: q = 35;
      432, 433, 434, 435, 436, 437, 438, 439, 440, 441, 442, 443: q = 36;
      444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455: q = 37;
      456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467: q = 38;
      468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479: q = 39;
      480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491: q = 40;
      492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503: q = 41;
      504, 505, 506, 507, 508, 509, 510, 511, 512, 513, 514, 515: q = 42;
      516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527: q = 43;
      528, 529, 530, 531, 532, 533, 534, 535, 536, 537, 538, 539: q = 44;
      540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551: q = 45;
      552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563: q = 46;
      564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575: q = 47;
      576, 577, 578, 579, 580, 581, 582, 583, 584, 585, 586, 587: q = 48;
      588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599: q = 49;
      600, 601, 602, 603, 604, 605, 606, 607, 608, 609, 610, 611: q = 50;
      612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 623: q = 51;
      624, 625, 626, 627, 628, 629, 630, 631, 632, 633, 634, 635: q = 52;
      636, 637, 638, 639, 640, 641, 642, 643, 644, 645, 646, 647: q = 53;
      648, 649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659: q = 54;
      660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670, 671: q = 55;
      672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683: q = 56;
      684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 695: q = 57;
      696, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707: q = 58;
      708, 709, 710, 711, 712, 713, 714, 715, 716, 717, 718, 719: q = 59;
      720, 721, 722, 723, 724, 725, 726, 727, 728, 729, 730, 731: q = 60;
      732, 733, 734, 735, 736, 737, 738, 739, 740, 741, 742, 743: q = 61;
      744, 745, 746, 747, 748, 749, 750, 751, 752, 753, 754, 755: q = 62;
      756, 757, 758, 759, 760, 761, 762, 763, 764, 765, 766, 767: q = 63;
      768, 769, 770, 771, 772, 773, 774, 775, 776, 777, 778, 779: q = 64;
      780, 781, 782, 783, 784, 785, 786, 787, 788, 789, 790, 791: q = 65;
      792, 793, 794, 795, 796, 797, 798, 799, 800, 801, 802, 803: q = 66;
      804, 805, 806, 807, 808, 809, 810, 811, 812, 813, 814, 815: q = 67;
      816, 817, 818, 819, 820, 821, 822, 823, 824, 825, 826, 827: q = 68;
      828, 829, 830, 831, 832, 833, 834, 835, 836, 837, 838, 839: q = 69;
      840, 841, 842, 843, 844, 845, 846, 847, 848, 849, 850, 851: q = 70;
      852, 853, 854, 855, 856, 857, 858, 859, 860, 861, 862, 863: q = 71;
      864, 865, 866, 867, 868, 869, 870, 871, 872, 873, 874, 875: q = 72;
      876, 877, 878, 879, 880, 881, 882, 883, 884, 885, 886, 887: q = 73;
      888, 889, 890, 891, 892, 893, 894, 895, 896, 897, 898, 899: q = 74;
      900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911: q = 75;
      912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923: q = 76;
      924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935: q = 77;
      936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947: q = 78;
      948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959: q = 79;
      960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971: q = 80;
      972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983: q = 81;
      984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995: q = 82;
      996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007:
      q = 83;
      1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019:
      q = 84;
      1020, 1021, 1022, 1023: q = 85;
      default: q = 8'dx;
    endcase
  end
endmodule