module CC (
  input clk,
  input rst_n,
  input in_valid,
  input [1:0] mode,
  input signed [7:0] xi,  // -128~127
  input signed [7:0] yi,  // -128~127
  output reg out_valid,
  output reg signed [7:0] xo,
  output reg signed [7:0] yo
);

  reg [2:0] state;
  localparam IDEL = 0, EAT = 1, OUT_mode0 = 2, PREOUT_1 = 3, PREOUT_2=4, OUT_mode1=5, OUT_mode2=6;

  reg [1:0] EATcnt;
  reg signed [7:0] p[0:3][1:2];
  reg signed [12:0] _reg[1:4];  // 13位
  reg signed [8:0] mul1[1:2];  // mode1, 2只要8位元, 0要9位元
  reg signed [8:0] mul2[1:2];  // mode1要14位
  wire signed [16:0] prod1 = mul1[1] * mul1[2];  // mode0要17位
  wire signed [16:0] prod2 = mul2[1] * mul2[2];  // mode0要17位
  wire cmp = _reg[1] < _reg[2];
  //************** for mode0 **************************
  reg signed [7:0] head, pos_x;
  reg signed [8:0] y_diff;  // 9位
  wire signed [8:0] a1_minus_c1 = p[0][1] - p[2][1];
  wire signed [8:0] a2_minus_c2 = p[0][2] - p[2][2];
  wire cmp_prod12 = prod1 > prod2;
  reg signed [8:0] r;  // 9位
  reg signed [7:0] offset;  // 8位
  wire signed [9:0] r_plus = r + a1_minus_c1;  // 10位
  wire signed [2:0] quotient = r_plus / a2_minus_c2;  // 3位
  wire signed [8:0] remainder = r_plus % a2_minus_c2;  // 9位

  // integer i;
  // reg [9:0] quotient;
  // reg [8:0] remainder;
  // reg [18:0] dividend, divisor;  // 10位除以9位
  // always @(*) begin
  //   dividend = r_plus;
  //   divisor  = {a2_minus_c2, 10'd0};
  //   for (i = 0; i < 10; i = i + 1) begin
  //     dividend = (dividend << 1);
  //     if (dividend[18:10] >= a2_minus_c2)
  //       dividend = dividend - divisor + 1;
  //   end
  //   quotient  = dividend[2:0];
  //   remainder = dividend[18:10];
  // end
  //************** for mode1 **************************
  wire [6:0] root;
  wire signed [5:0] signx = xi[5:0];
  wire signed [5:0] signy = yi[5:0];
  wire signed [5:0] a2_minus_b2 = $signed(p[0][2][5:0]) - signy;
  wire signed [5:0] b1_minus_a1 = signx - $signed(p[0][1][5:0]);
  wire signed [16:0] prod1_minus_prod2 = prod1 - prod2;// 原始25位 mode2只要16位
  //************** for mode2 ************************
  reg signed [16:0] area;
  wire signed [16:0] area_next = area + prod1_minus_prod2;
  wire lastpoint = (xo == p[1][1] && yo == p[1][2]);

  // Mode0: Trapezoid rendering 
  //  輸入依序為 左上、右上、左下、右下，輸出要從左到右，最下排先
  //  只要方格有任一點被嚴格包在梯形內部就算，並且剛好只削到格子左下的話也算包到(此狀況只會出現在上邊跟右邊)
  //  定義線段ab，則點p與ab之間的關係為：
  //  (b1-a1)(p1-a2) > (b2-a2)(p0-a1) => 點在左邊
  //  (b1-a1)(p1-a2) > (b2-a2)(p0-a1) => 點在右邊
  //  (b1-a1)(p1-a2) = (b2-a2)(p0-a1) => 點在線上
  //  pattern 在 input.txt & ans.txt
  // Mode1: Relationship of a circle and a line
  //  輸入依序為直線端點a、直線端點b、圓心c、圓邊d，座標都是6bit二補數 -32 ~ 31
  //  要判斷[(a2-b2)c1 + (b1-a1)c2 + (a1b2-a2b1)]^2 與
  //  [(d1-c1)^2 + (d2-c2)^2][(a2-b2)^2 + (b1-a1)^2]的關係
  //  前者是距離平方，後者是半徑平方(<=7938^2)，是個平方VS積的問題
  //  外離{xo,yo}={0,0}，內割{xo,yo}={0,1}，相切{xo,yo}={0,2}
  //  b出:a2-b2, b1-a1, a1b2-a2b1,  (a2-b2)^2, (b1-a1)^2
  //  c出:(a2-b2)c1+(b1-a1)c2及大平方[.. + (a1b2-a2b1)]^2
  //  d出:(d1-c1)^2 (d2-c2)^2及[12位]*[12位]  2個小平方器及24位cmp
  //  pattern 在 coordinate_in.txt & coordinate_out.txt

  // r
  always @(posedge clk) begin
    if (EATcnt == 3) r <= 0;
    else if ((state == OUT_mode0 && !out_valid) || cmp_prod12) r <= remainder;
  end
  // offset
  always @(posedge clk) begin
    if (EATcnt == 3) offset <= 0;
    else if ((state == OUT_mode0 && !out_valid) || cmp_prod12)
      offset <= offset + quotient;
  end
  // head
  always @(*) begin
    head = r < 0 ? p[2][1] + offset - 1 : p[2][1] + offset;
  end
  // pos_x
  always @(posedge clk) begin
    if (state == OUT_mode0 && !out_valid) pos_x <= p[2][1];  // c1
    else if (cmp_prod12)  //(x-d1)(b2-d2) > (b1-d1)*y_diff列尾失效
      pos_x <= head;
    else  // (x-d1)(b2-d2)<=(b1-d1)(y_diff-1)列尾ok
      pos_x <= pos_x + 1;
  end
  // y_diff
  always @(posedge clk) begin
    if (EATcnt == 3) y_diff <= 1;
    else if (state==OUT_mode0 && out_valid && cmp_prod12) //(x-d1)(b2-d2) > (b1-d1)*y_diff列尾失效 
      y_diff <= y_diff + 1;
  end

  wire [5:0] abs_a2b2 = _reg[1][12] ? (~_reg[1]) + 6'd1 : _reg[1];
  wire [5:0] abs_b1a1 = _reg[2][12] ? (~_reg[2]) + 6'd1 : _reg[2];
  wire [5:0] ab_smaller = abs_b1a1 > abs_a2b2 ? abs_a2b2 : abs_b1a1;
  wire [5:0] ab_larger = abs_a2b2 > abs_b1a1 ? abs_a2b2 : abs_b1a1;

  wire [5:0] abs_d1c1 = p[3][1] > p[2][1] ? p[3][1] - p[2][1] : p[2][1] - p[3][1];
  wire [5:0] abs_d2c2 = p[3][2] > p[2][2] ? p[3][2] - p[2][2] : p[2][2] - p[3][2];
  wire [5:0] cd_smaller = abs_d1c1 > abs_d2c2 ? abs_d2c2 : abs_d1c1;
  wire [5:0] cd_larger = abs_d1c1 > abs_d2c2 ? abs_d1c1 : abs_d2c2;

  wire [5:0] smaller = EATcnt[1] ^ EATcnt[0] ? ab_smaller : cd_smaller;
  wire [5:0] larger = EATcnt[1] ^ EATcnt[0] ? ab_larger : cd_larger;

  root_module ABCD (
    smaller,
    larger,
    root
  );

  // _reg
  always @(posedge clk) begin
    if ((state == EAT) || state == PREOUT_1) begin
      if (EATcnt == 0) begin  // 輸出
        _reg[1] <= _reg[1][12] ? (~_reg[1]) + 13'd1 : _reg[1];
        _reg[2] <= prod2;  // root_ab * root_cd
        // _reg[2] <= _reg[4] * root;  // root_ab * root_cd
      end else if (EATcnt == 3) begin  // 正d
        _reg[1] <= $signed(
          _reg[1][11:0]
        ) + $signed(
          _reg[2][11:0]
        ) + $signed(
          _reg[3][11:0]
        );  // (a2-b2)c1 + (b1-a1)c2 + (a1b2-a2b1)
        // _reg[3] <= root;  // root_cd
      end else if (EATcnt == 2) begin  // 正c
        _reg[1] <= prod1;  // (a2-b2)c1
        _reg[2] <= prod2;  // (b1-a1)c2
        _reg[4] <= root;  // root_ab 45
      end else if (EATcnt == 1) begin  // 正b
        _reg[1] <= p[0][2] - yi;  // a2-b2
        _reg[2] <= xi - p[0][1];  // b1-a1
        _reg[3] <= prod1_minus_prod2;  //a1b2-a2b1
      end
    end
  end
  // mul1
  always @(*) begin
    if (state == OUT_mode0) begin
      mul1[1] = pos_x + 1 - p[3][1];  // x - d1
      mul1[2] = p[1][2] - p[3][2];  // (b2-d2)
    end else if (state == EAT && mode == 1) begin
      if (EATcnt == 1) begin  // 吃b前
        mul1[1] = p[0][1];  // a1
        mul1[2] = signy;  // b2
      end else if (EATcnt == 2) begin  // 吃c前
        mul1[1] = _reg[1];  // (a2-b2)
        mul1[2] = signx;  // c1
      end else begin
        mul1[1] = 9'dx;
        mul1[2] = 9'dx;
      end
    end else if (state == PREOUT_2) begin
      mul1[1] = p[3][1];  // d1
      mul1[2] = p[0][2];  // a2
    end else if (state == EAT && mode == 2) begin
      mul1[1] = p[EATcnt-1][1];
      mul1[2] = yi;
    end else begin
      mul1[1] = 9'dx;
      mul1[2] = 9'dx;
    end
  end

  // mul2
  always @(*) begin
    if (state == PREOUT_2) begin
      mul2[1] = p[3][2];  // d2
      mul2[2] = p[0][1];  // a1
    end else if (state == OUT_mode0) begin
      mul2[1] = p[1][1] - p[3][1];  // b1-d1
      mul2[2] = y_diff - 1;  // y_diff_now
    end else if ((mode == 1) || state == PREOUT_1) begin
      if (EATcnt == 2) begin  // 吃c前
        mul2[1] = _reg[2];  // b1-a1
        mul2[2] = signy;  // c2
      end else if (EATcnt == 1) begin  // 吃b前
        mul2[1] = p[0][2];  // a2
        mul2[2] = signx;  // b1
      end else begin
        mul2[1] = _reg[4];  // root_ab
        mul2[2] = root;  // root_cd
      end
    end else if (state == EAT && mode == 2) begin
      mul2[1] = p[EATcnt-1][2];
      mul2[2] = xi;
    end else begin
      mul2[1] = 9'dx;
      mul2[2] = 9'dx;
    end
  end

  // p[i][1], p[i][2]
  always @(posedge clk) begin
    if (in_valid) {p[EATcnt][1], p[EATcnt][2]} <= {xi, yi};
  end
  // EATcnt 0吃a  1吃b  2吃c  3吃d
  always @(posedge clk, negedge rst_n) begin
    if (!rst_n) EATcnt <= 0;
    else if (in_valid) EATcnt <= EATcnt + 1;
  end

  // area
  always @(posedge clk, negedge rst_n) begin
    if (!rst_n) area <= 0;
    else if (state == PREOUT_2)
      area <= (area_next[16]) ?  // 負的面積
      (~(area_next) + 1) >> 1 : (area_next) >> 1;
    else if (state == EAT) begin
      area <= area_next;
    end else area <= 0;
  end

  // xo, yo
  always @(*) begin
    if (state == OUT_mode1) begin
      xo = 0;
      yo = {6'd0, _reg[1] == _reg[2], cmp};
    end else if (state == OUT_mode0) begin
      xo = pos_x;
      yo = p[2][2] + y_diff - 1;
    end else if (state == OUT_mode2) begin
      {xo, yo} = area;
    end else begin
      {xo, yo} = 0;
    end
  end

  // state
  always @(posedge clk, negedge rst_n) begin
    if (!rst_n) state <= IDEL;
    else if (state == OUT_mode0 && !lastpoint) state <= OUT_mode0;
    else if (EATcnt == 3) begin  // 正d
      case (mode)
        0: state <= OUT_mode0;
        1: state <= PREOUT_1;
        2: state <= PREOUT_2;
      endcase
    end else if (in_valid) state <= EAT;
    else begin
      case (state)
        PREOUT_1: state <= OUT_mode1;
        PREOUT_2: state <= OUT_mode2;
        default:  state <= IDEL;
      endcase
    end
  end


  // out_valid
  always @(posedge clk, negedge rst_n) begin
    if (!rst_n) out_valid <= 0;
    else if ((state == OUT_mode0 && !lastpoint) 
    || state == PREOUT_1
    || state == PREOUT_2)
      out_valid <= 1'b1;
    else out_valid <= 0;
  end
  // Mode2: Calculate the area of a quadrilateral
  //  順時鐘依序輸入點a、點b、點c、點d
  //  面積=(1/2)*[(a1b2-a2b1)+(b1c2-b2c1)+(c1d2-c2d1)+(d1a2-d2a1)]向下取整
  //  pattern 在 area_in.txt & area_out.txt

endmodule

module root_module (
  input [5:0] a,
  input [5:0] b,
  output reg [6:0] c
);

  // always @(*) begin
  //   c = b + ((3 * a) >> 3);
  // end
  always @(*) begin
    case ({
      a, b
    })
      {6'd0, 6'd0} : c = 0;
      {6'd0, 6'd1} : c = 1;
      {6'd0, 6'd2} : c = 2;
      {6'd0, 6'd3} : c = 3;
      {6'd0, 6'd4} : c = 4;
      {6'd0, 6'd5} : c = 5;
      {6'd0, 6'd6} : c = 6;
      {6'd0, 6'd7} : c = 7;
      {6'd0, 6'd8} : c = 8;
      {6'd0, 6'd9} : c = 9;
      {6'd0, 6'd10} : c = 10;
      {6'd0, 6'd11} : c = 11;
      {6'd0, 6'd12} : c = 12;
      {6'd0, 6'd13} : c = 13;
      {6'd0, 6'd14} : c = 14;
      {6'd0, 6'd15} : c = 15;
      {6'd0, 6'd16} : c = 16;
      {6'd0, 6'd17} : c = 17;
      {6'd0, 6'd18} : c = 18;
      {6'd0, 6'd19} : c = 19;
      {6'd0, 6'd20} : c = 20;
      {6'd0, 6'd21} : c = 21;
      {6'd0, 6'd22} : c = 22;
      {6'd0, 6'd23} : c = 23;
      {6'd0, 6'd24} : c = 24;
      {6'd0, 6'd25} : c = 25;
      {6'd0, 6'd26} : c = 26;
      {6'd0, 6'd27} : c = 27;
      {6'd0, 6'd28} : c = 28;
      {6'd0, 6'd29} : c = 29;
      {6'd0, 6'd30} : c = 30;
      {6'd0, 6'd31} : c = 31;
      {6'd0, 6'd32} : c = 32;
      {6'd0, 6'd33} : c = 33;
      {6'd0, 6'd34} : c = 34;
      {6'd0, 6'd35} : c = 35;
      {6'd0, 6'd36} : c = 36;
      {6'd0, 6'd37} : c = 37;
      {6'd0, 6'd38} : c = 38;
      {6'd0, 6'd39} : c = 39;
      {6'd0, 6'd40} : c = 40;
      {6'd0, 6'd41} : c = 41;
      {6'd0, 6'd42} : c = 42;
      {6'd0, 6'd43} : c = 43;
      {6'd0, 6'd44} : c = 44;
      {6'd0, 6'd45} : c = 45;
      {6'd0, 6'd46} : c = 46;
      {6'd0, 6'd47} : c = 47;
      {6'd0, 6'd48} : c = 48;
      {6'd0, 6'd49} : c = 49;
      {6'd0, 6'd50} : c = 50;
      {6'd0, 6'd51} : c = 51;
      {6'd0, 6'd52} : c = 52;
      {6'd0, 6'd53} : c = 53;
      {6'd0, 6'd54} : c = 54;
      {6'd0, 6'd55} : c = 55;
      {6'd0, 6'd56} : c = 56;
      {6'd0, 6'd57} : c = 57;
      {6'd0, 6'd58} : c = 58;
      {6'd0, 6'd59} : c = 59;
      {6'd0, 6'd60} : c = 60;
      {6'd0, 6'd61} : c = 61;
      {6'd0, 6'd62} : c = 62;
      {6'd0, 6'd63} : c = 63;
      {6'd1, 6'd1} : c = 1;
      {6'd1, 6'd2} : c = 2;
      {6'd1, 6'd3} : c = 3;
      {6'd1, 6'd4} : c = 4;
      {6'd1, 6'd5} : c = 5;
      {6'd1, 6'd6} : c = 6;
      {6'd1, 6'd7} : c = 7;
      {6'd1, 6'd8} : c = 8;
      {6'd1, 6'd9} : c = 9;
      {6'd1, 6'd10} : c = 10;
      {6'd1, 6'd11} : c = 11;
      {6'd1, 6'd12} : c = 12;
      {6'd1, 6'd13} : c = 13;
      {6'd1, 6'd14} : c = 14;
      {6'd1, 6'd15} : c = 15;
      {6'd1, 6'd16} : c = 16;
      {6'd1, 6'd17} : c = 17;
      {6'd1, 6'd18} : c = 18;
      {6'd1, 6'd19} : c = 19;
      {6'd1, 6'd20} : c = 20;
      {6'd1, 6'd21} : c = 21;
      {6'd1, 6'd22} : c = 22;
      {6'd1, 6'd23} : c = 23;
      {6'd1, 6'd24} : c = 24;
      {6'd1, 6'd25} : c = 25;
      {6'd1, 6'd26} : c = 26;
      {6'd1, 6'd27} : c = 27;
      {6'd1, 6'd28} : c = 28;
      {6'd1, 6'd29} : c = 29;
      {6'd1, 6'd30} : c = 30;
      {6'd1, 6'd31} : c = 31;
      {6'd1, 6'd32} : c = 32;
      {6'd1, 6'd33} : c = 33;
      {6'd1, 6'd34} : c = 34;
      {6'd1, 6'd35} : c = 35;
      {6'd1, 6'd36} : c = 36;
      {6'd1, 6'd37} : c = 37;
      {6'd1, 6'd38} : c = 38;
      {6'd1, 6'd39} : c = 39;
      {6'd1, 6'd40} : c = 40;
      {6'd1, 6'd41} : c = 41;
      {6'd1, 6'd42} : c = 42;
      {6'd1, 6'd43} : c = 43;
      {6'd1, 6'd44} : c = 44;
      {6'd1, 6'd45} : c = 45;
      {6'd1, 6'd46} : c = 46;
      {6'd1, 6'd47} : c = 47;
      {6'd1, 6'd48} : c = 48;
      {6'd1, 6'd49} : c = 49;
      {6'd1, 6'd50} : c = 50;
      {6'd1, 6'd51} : c = 51;
      {6'd1, 6'd52} : c = 52;
      {6'd1, 6'd53} : c = 53;
      {6'd1, 6'd54} : c = 54;
      {6'd1, 6'd55} : c = 55;
      {6'd1, 6'd56} : c = 56;
      {6'd1, 6'd57} : c = 57;
      {6'd1, 6'd58} : c = 58;
      {6'd1, 6'd59} : c = 59;
      {6'd1, 6'd60} : c = 60;
      {6'd1, 6'd61} : c = 61;
      {6'd1, 6'd62} : c = 62;
      {6'd1, 6'd63} : c = 63;
      {6'd2, 6'd2} : c = 3;
      {6'd2, 6'd3} : c = 4;
      {6'd2, 6'd4} : c = 4;
      {6'd2, 6'd5} : c = 5;
      {6'd2, 6'd6} : c = 6;
      {6'd2, 6'd7} : c = 7;
      {6'd2, 6'd8} : c = 8;
      {6'd2, 6'd9} : c = 9;
      {6'd2, 6'd10} : c = 10;
      {6'd2, 6'd11} : c = 11;
      {6'd2, 6'd12} : c = 12;
      {6'd2, 6'd13} : c = 13;
      {6'd2, 6'd14} : c = 14;
      {6'd2, 6'd15} : c = 15;
      {6'd2, 6'd16} : c = 16;
      {6'd2, 6'd17} : c = 17;
      {6'd2, 6'd18} : c = 18;
      {6'd2, 6'd19} : c = 19;
      {6'd2, 6'd20} : c = 20;
      {6'd2, 6'd21} : c = 21;
      {6'd2, 6'd22} : c = 22;
      {6'd2, 6'd23} : c = 23;
      {6'd2, 6'd24} : c = 24;
      {6'd2, 6'd25} : c = 25;
      {6'd2, 6'd26} : c = 26;
      {6'd2, 6'd27} : c = 27;
      {6'd2, 6'd28} : c = 28;
      {6'd2, 6'd29} : c = 29;
      {6'd2, 6'd30} : c = 30;
      {6'd2, 6'd31} : c = 31;
      {6'd2, 6'd32} : c = 32;
      {6'd2, 6'd33} : c = 33;
      {6'd2, 6'd34} : c = 34;
      {6'd2, 6'd35} : c = 35;
      {6'd2, 6'd36} : c = 36;
      {6'd2, 6'd37} : c = 37;
      {6'd2, 6'd38} : c = 38;
      {6'd2, 6'd39} : c = 39;
      {6'd2, 6'd40} : c = 40;
      {6'd2, 6'd41} : c = 41;
      {6'd2, 6'd42} : c = 42;
      {6'd2, 6'd43} : c = 43;
      {6'd2, 6'd44} : c = 44;
      {6'd2, 6'd45} : c = 45;
      {6'd2, 6'd46} : c = 46;
      {6'd2, 6'd47} : c = 47;
      {6'd2, 6'd48} : c = 48;
      {6'd2, 6'd49} : c = 49;
      {6'd2, 6'd50} : c = 50;
      {6'd2, 6'd51} : c = 51;
      {6'd2, 6'd52} : c = 52;
      {6'd2, 6'd53} : c = 53;
      {6'd2, 6'd54} : c = 54;
      {6'd2, 6'd55} : c = 55;
      {6'd2, 6'd56} : c = 56;
      {6'd2, 6'd57} : c = 57;
      {6'd2, 6'd58} : c = 58;
      {6'd2, 6'd59} : c = 59;
      {6'd2, 6'd60} : c = 60;
      {6'd2, 6'd61} : c = 61;
      {6'd2, 6'd62} : c = 62;
      {6'd2, 6'd63} : c = 63;
      {6'd3, 6'd3} : c = 4;
      {6'd3, 6'd4} : c = 5;
      {6'd3, 6'd5} : c = 6;
      {6'd3, 6'd6} : c = 7;
      {6'd3, 6'd7} : c = 8;
      {6'd3, 6'd8} : c = 9;
      {6'd3, 6'd9} : c = 9;
      {6'd3, 6'd10} : c = 10;
      {6'd3, 6'd11} : c = 11;
      {6'd3, 6'd12} : c = 12;
      {6'd3, 6'd13} : c = 13;
      {6'd3, 6'd14} : c = 14;
      {6'd3, 6'd15} : c = 15;
      {6'd3, 6'd16} : c = 16;
      {6'd3, 6'd17} : c = 17;
      {6'd3, 6'd18} : c = 18;
      {6'd3, 6'd19} : c = 19;
      {6'd3, 6'd20} : c = 20;
      {6'd3, 6'd21} : c = 21;
      {6'd3, 6'd22} : c = 22;
      {6'd3, 6'd23} : c = 23;
      {6'd3, 6'd24} : c = 24;
      {6'd3, 6'd25} : c = 25;
      {6'd3, 6'd26} : c = 26;
      {6'd3, 6'd27} : c = 27;
      {6'd3, 6'd28} : c = 28;
      {6'd3, 6'd29} : c = 29;
      {6'd3, 6'd30} : c = 30;
      {6'd3, 6'd31} : c = 31;
      {6'd3, 6'd32} : c = 32;
      {6'd3, 6'd33} : c = 33;
      {6'd3, 6'd34} : c = 34;
      {6'd3, 6'd35} : c = 35;
      {6'd3, 6'd36} : c = 36;
      {6'd3, 6'd37} : c = 37;
      {6'd3, 6'd38} : c = 38;
      {6'd3, 6'd39} : c = 39;
      {6'd3, 6'd40} : c = 40;
      {6'd3, 6'd41} : c = 41;
      {6'd3, 6'd42} : c = 42;
      {6'd3, 6'd43} : c = 43;
      {6'd3, 6'd44} : c = 44;
      {6'd3, 6'd45} : c = 45;
      {6'd3, 6'd46} : c = 46;
      {6'd3, 6'd47} : c = 47;
      {6'd3, 6'd48} : c = 48;
      {6'd3, 6'd49} : c = 49;
      {6'd3, 6'd50} : c = 50;
      {6'd3, 6'd51} : c = 51;
      {6'd3, 6'd52} : c = 52;
      {6'd3, 6'd53} : c = 53;
      {6'd3, 6'd54} : c = 54;
      {6'd3, 6'd55} : c = 55;
      {6'd3, 6'd56} : c = 56;
      {6'd3, 6'd57} : c = 57;
      {6'd3, 6'd58} : c = 58;
      {6'd3, 6'd59} : c = 59;
      {6'd3, 6'd60} : c = 60;
      {6'd3, 6'd61} : c = 61;
      {6'd3, 6'd62} : c = 62;
      {6'd3, 6'd63} : c = 63;
      {6'd4, 6'd4} : c = 6;
      {6'd4, 6'd5} : c = 6;
      {6'd4, 6'd6} : c = 7;
      {6'd4, 6'd7} : c = 8;
      {6'd4, 6'd8} : c = 9;
      {6'd4, 6'd9} : c = 10;
      {6'd4, 6'd10} : c = 11;
      {6'd4, 6'd11} : c = 12;
      {6'd4, 6'd12} : c = 13;
      {6'd4, 6'd13} : c = 14;
      {6'd4, 6'd14} : c = 15;
      {6'd4, 6'd15} : c = 16;
      {6'd4, 6'd16} : c = 16;
      {6'd4, 6'd17} : c = 17;
      {6'd4, 6'd18} : c = 18;
      {6'd4, 6'd19} : c = 19;
      {6'd4, 6'd20} : c = 20;
      {6'd4, 6'd21} : c = 21;
      {6'd4, 6'd22} : c = 22;
      {6'd4, 6'd23} : c = 23;
      {6'd4, 6'd24} : c = 24;
      {6'd4, 6'd25} : c = 25;
      {6'd4, 6'd26} : c = 26;
      {6'd4, 6'd27} : c = 27;
      {6'd4, 6'd28} : c = 28;
      {6'd4, 6'd29} : c = 29;
      {6'd4, 6'd30} : c = 30;
      {6'd4, 6'd31} : c = 31;
      {6'd4, 6'd32} : c = 32;
      {6'd4, 6'd33} : c = 33;
      {6'd4, 6'd34} : c = 34;
      {6'd4, 6'd35} : c = 35;
      {6'd4, 6'd36} : c = 36;
      {6'd4, 6'd37} : c = 37;
      {6'd4, 6'd38} : c = 38;
      {6'd4, 6'd39} : c = 39;
      {6'd4, 6'd40} : c = 40;
      {6'd4, 6'd41} : c = 41;
      {6'd4, 6'd42} : c = 42;
      {6'd4, 6'd43} : c = 43;
      {6'd4, 6'd44} : c = 44;
      {6'd4, 6'd45} : c = 45;
      {6'd4, 6'd46} : c = 46;
      {6'd4, 6'd47} : c = 47;
      {6'd4, 6'd48} : c = 48;
      {6'd4, 6'd49} : c = 49;
      {6'd4, 6'd50} : c = 50;
      {6'd4, 6'd51} : c = 51;
      {6'd4, 6'd52} : c = 52;
      {6'd4, 6'd53} : c = 53;
      {6'd4, 6'd54} : c = 54;
      {6'd4, 6'd55} : c = 55;
      {6'd4, 6'd56} : c = 56;
      {6'd4, 6'd57} : c = 57;
      {6'd4, 6'd58} : c = 58;
      {6'd4, 6'd59} : c = 59;
      {6'd4, 6'd60} : c = 60;
      {6'd4, 6'd61} : c = 61;
      {6'd4, 6'd62} : c = 62;
      {6'd4, 6'd63} : c = 63;
      {6'd5, 6'd5} : c = 7;
      {6'd5, 6'd6} : c = 8;
      {6'd5, 6'd7} : c = 9;
      {6'd5, 6'd8} : c = 9;
      {6'd5, 6'd9} : c = 10;
      {6'd5, 6'd10} : c = 11;
      {6'd5, 6'd11} : c = 12;
      {6'd5, 6'd12} : c = 13;
      {6'd5, 6'd13} : c = 14;
      {6'd5, 6'd14} : c = 15;
      {6'd5, 6'd15} : c = 16;
      {6'd5, 6'd16} : c = 17;
      {6'd5, 6'd17} : c = 18;
      {6'd5, 6'd18} : c = 19;
      {6'd5, 6'd19} : c = 20;
      {6'd5, 6'd20} : c = 21;
      {6'd5, 6'd21} : c = 22;
      {6'd5, 6'd22} : c = 23;
      {6'd5, 6'd23} : c = 24;
      {6'd5, 6'd24} : c = 25;
      {6'd5, 6'd25} : c = 25;
      {6'd5, 6'd26} : c = 26;
      {6'd5, 6'd27} : c = 27;
      {6'd5, 6'd28} : c = 28;
      {6'd5, 6'd29} : c = 29;
      {6'd5, 6'd30} : c = 30;
      {6'd5, 6'd31} : c = 31;
      {6'd5, 6'd32} : c = 32;
      {6'd5, 6'd33} : c = 33;
      {6'd5, 6'd34} : c = 34;
      {6'd5, 6'd35} : c = 35;
      {6'd5, 6'd36} : c = 36;
      {6'd5, 6'd37} : c = 37;
      {6'd5, 6'd38} : c = 38;
      {6'd5, 6'd39} : c = 39;
      {6'd5, 6'd40} : c = 40;
      {6'd5, 6'd41} : c = 41;
      {6'd5, 6'd42} : c = 42;
      {6'd5, 6'd43} : c = 43;
      {6'd5, 6'd44} : c = 44;
      {6'd5, 6'd45} : c = 45;
      {6'd5, 6'd46} : c = 46;
      {6'd5, 6'd47} : c = 47;
      {6'd5, 6'd48} : c = 48;
      {6'd5, 6'd49} : c = 49;
      {6'd5, 6'd50} : c = 50;
      {6'd5, 6'd51} : c = 51;
      {6'd5, 6'd52} : c = 52;
      {6'd5, 6'd53} : c = 53;
      {6'd5, 6'd54} : c = 54;
      {6'd5, 6'd55} : c = 55;
      {6'd5, 6'd56} : c = 56;
      {6'd5, 6'd57} : c = 57;
      {6'd5, 6'd58} : c = 58;
      {6'd5, 6'd59} : c = 59;
      {6'd5, 6'd60} : c = 60;
      {6'd5, 6'd61} : c = 61;
      {6'd5, 6'd62} : c = 62;
      {6'd5, 6'd63} : c = 63;
      {6'd6, 6'd6} : c = 8;
      {6'd6, 6'd7} : c = 9;
      {6'd6, 6'd8} : c = 10;
      {6'd6, 6'd9} : c = 11;
      {6'd6, 6'd10} : c = 12;
      {6'd6, 6'd11} : c = 13;
      {6'd6, 6'd12} : c = 13;
      {6'd6, 6'd13} : c = 14;
      {6'd6, 6'd14} : c = 15;
      {6'd6, 6'd15} : c = 16;
      {6'd6, 6'd16} : c = 17;
      {6'd6, 6'd17} : c = 18;
      {6'd6, 6'd18} : c = 19;
      {6'd6, 6'd19} : c = 20;
      {6'd6, 6'd20} : c = 21;
      {6'd6, 6'd21} : c = 22;
      {6'd6, 6'd22} : c = 23;
      {6'd6, 6'd23} : c = 24;
      {6'd6, 6'd24} : c = 25;
      {6'd6, 6'd25} : c = 26;
      {6'd6, 6'd26} : c = 27;
      {6'd6, 6'd27} : c = 28;
      {6'd6, 6'd28} : c = 29;
      {6'd6, 6'd29} : c = 30;
      {6'd6, 6'd30} : c = 31;
      {6'd6, 6'd31} : c = 32;
      {6'd6, 6'd32} : c = 33;
      {6'd6, 6'd33} : c = 34;
      {6'd6, 6'd34} : c = 35;
      {6'd6, 6'd35} : c = 36;
      {6'd6, 6'd36} : c = 36;
      {6'd6, 6'd37} : c = 37;
      {6'd6, 6'd38} : c = 38;
      {6'd6, 6'd39} : c = 39;
      {6'd6, 6'd40} : c = 40;
      {6'd6, 6'd41} : c = 41;
      {6'd6, 6'd42} : c = 42;
      {6'd6, 6'd43} : c = 43;
      {6'd6, 6'd44} : c = 44;
      {6'd6, 6'd45} : c = 45;
      {6'd6, 6'd46} : c = 46;
      {6'd6, 6'd47} : c = 47;
      {6'd6, 6'd48} : c = 48;
      {6'd6, 6'd49} : c = 49;
      {6'd6, 6'd50} : c = 50;
      {6'd6, 6'd51} : c = 51;
      {6'd6, 6'd52} : c = 52;
      {6'd6, 6'd53} : c = 53;
      {6'd6, 6'd54} : c = 54;
      {6'd6, 6'd55} : c = 55;
      {6'd6, 6'd56} : c = 56;
      {6'd6, 6'd57} : c = 57;
      {6'd6, 6'd58} : c = 58;
      {6'd6, 6'd59} : c = 59;
      {6'd6, 6'd60} : c = 60;
      {6'd6, 6'd61} : c = 61;
      {6'd6, 6'd62} : c = 62;
      {6'd6, 6'd63} : c = 63;
      {6'd7, 6'd7} : c = 10;
      {6'd7, 6'd8} : c = 11;
      {6'd7, 6'd9} : c = 11;
      {6'd7, 6'd10} : c = 12;
      {6'd7, 6'd11} : c = 13;
      {6'd7, 6'd12} : c = 14;
      {6'd7, 6'd13} : c = 15;
      {6'd7, 6'd14} : c = 16;
      {6'd7, 6'd15} : c = 17;
      {6'd7, 6'd16} : c = 17;
      {6'd7, 6'd17} : c = 18;
      {6'd7, 6'd18} : c = 19;
      {6'd7, 6'd19} : c = 20;
      {6'd7, 6'd20} : c = 21;
      {6'd7, 6'd21} : c = 22;
      {6'd7, 6'd22} : c = 23;
      {6'd7, 6'd23} : c = 24;
      {6'd7, 6'd24} : c = 25;
      {6'd7, 6'd25} : c = 26;
      {6'd7, 6'd26} : c = 27;
      {6'd7, 6'd27} : c = 28;
      {6'd7, 6'd28} : c = 29;
      {6'd7, 6'd29} : c = 30;
      {6'd7, 6'd30} : c = 31;
      {6'd7, 6'd31} : c = 32;
      {6'd7, 6'd32} : c = 33;
      {6'd7, 6'd33} : c = 34;
      {6'd7, 6'd34} : c = 35;
      {6'd7, 6'd35} : c = 36;
      {6'd7, 6'd36} : c = 37;
      {6'd7, 6'd37} : c = 38;
      {6'd7, 6'd38} : c = 39;
      {6'd7, 6'd39} : c = 40;
      {6'd7, 6'd40} : c = 41;
      {6'd7, 6'd41} : c = 42;
      {6'd7, 6'd42} : c = 43;
      {6'd7, 6'd43} : c = 44;
      {6'd7, 6'd44} : c = 45;
      {6'd7, 6'd45} : c = 46;
      {6'd7, 6'd46} : c = 47;
      {6'd7, 6'd47} : c = 48;
      {6'd7, 6'd48} : c = 49;
      {6'd7, 6'd49} : c = 49;
      {6'd7, 6'd50} : c = 50;
      {6'd7, 6'd51} : c = 51;
      {6'd7, 6'd52} : c = 52;
      {6'd7, 6'd53} : c = 53;
      {6'd7, 6'd54} : c = 54;
      {6'd7, 6'd55} : c = 55;
      {6'd7, 6'd56} : c = 56;
      {6'd7, 6'd57} : c = 57;
      {6'd7, 6'd58} : c = 58;
      {6'd7, 6'd59} : c = 59;
      {6'd7, 6'd60} : c = 60;
      {6'd7, 6'd61} : c = 61;
      {6'd7, 6'd62} : c = 62;
      {6'd7, 6'd63} : c = 63;
      {6'd8, 6'd8} : c = 11;
      {6'd8, 6'd9} : c = 12;
      {6'd8, 6'd10} : c = 13;
      {6'd8, 6'd11} : c = 14;
      {6'd8, 6'd12} : c = 14;
      {6'd8, 6'd13} : c = 15;
      {6'd8, 6'd14} : c = 16;
      {6'd8, 6'd15} : c = 17;
      {6'd8, 6'd16} : c = 18;
      {6'd8, 6'd17} : c = 19;
      {6'd8, 6'd18} : c = 20;
      {6'd8, 6'd19} : c = 21;
      {6'd8, 6'd20} : c = 22;
      {6'd8, 6'd21} : c = 22;
      {6'd8, 6'd22} : c = 23;
      {6'd8, 6'd23} : c = 24;
      {6'd8, 6'd24} : c = 25;
      {6'd8, 6'd25} : c = 26;
      {6'd8, 6'd26} : c = 27;
      {6'd8, 6'd27} : c = 28;
      {6'd8, 6'd28} : c = 29;
      {6'd8, 6'd29} : c = 30;
      {6'd8, 6'd30} : c = 31;
      {6'd8, 6'd31} : c = 32;
      {6'd8, 6'd32} : c = 33;
      {6'd8, 6'd33} : c = 34;
      {6'd8, 6'd34} : c = 35;
      {6'd8, 6'd35} : c = 36;
      {6'd8, 6'd36} : c = 37;
      {6'd8, 6'd37} : c = 38;
      {6'd8, 6'd38} : c = 39;
      {6'd8, 6'd39} : c = 40;
      {6'd8, 6'd40} : c = 41;
      {6'd8, 6'd41} : c = 42;
      {6'd8, 6'd42} : c = 43;
      {6'd8, 6'd43} : c = 44;
      {6'd8, 6'd44} : c = 45;
      {6'd8, 6'd45} : c = 46;
      {6'd8, 6'd46} : c = 47;
      {6'd8, 6'd47} : c = 48;
      {6'd8, 6'd48} : c = 49;
      {6'd8, 6'd49} : c = 50;
      {6'd8, 6'd50} : c = 51;
      {6'd8, 6'd51} : c = 52;
      {6'd8, 6'd52} : c = 53;
      {6'd8, 6'd53} : c = 54;
      {6'd8, 6'd54} : c = 55;
      {6'd8, 6'd55} : c = 56;
      {6'd8, 6'd56} : c = 57;
      {6'd8, 6'd57} : c = 58;
      {6'd8, 6'd58} : c = 59;
      {6'd8, 6'd59} : c = 60;
      {6'd8, 6'd60} : c = 61;
      {6'd8, 6'd61} : c = 62;
      {6'd8, 6'd62} : c = 63;
      {6'd8, 6'd63} : c = 64;
      {6'd9, 6'd9} : c = 13;
      {6'd9, 6'd10} : c = 13;
      {6'd9, 6'd11} : c = 14;
      {6'd9, 6'd12} : c = 15;
      {6'd9, 6'd13} : c = 16;
      {6'd9, 6'd14} : c = 17;
      {6'd9, 6'd15} : c = 17;
      {6'd9, 6'd16} : c = 18;
      {6'd9, 6'd17} : c = 19;
      {6'd9, 6'd18} : c = 20;
      {6'd9, 6'd19} : c = 21;
      {6'd9, 6'd20} : c = 22;
      {6'd9, 6'd21} : c = 23;
      {6'd9, 6'd22} : c = 24;
      {6'd9, 6'd23} : c = 25;
      {6'd9, 6'd24} : c = 26;
      {6'd9, 6'd25} : c = 27;
      {6'd9, 6'd26} : c = 28;
      {6'd9, 6'd27} : c = 28;
      {6'd9, 6'd28} : c = 29;
      {6'd9, 6'd29} : c = 30;
      {6'd9, 6'd30} : c = 31;
      {6'd9, 6'd31} : c = 32;
      {6'd9, 6'd32} : c = 33;
      {6'd9, 6'd33} : c = 34;
      {6'd9, 6'd34} : c = 35;
      {6'd9, 6'd35} : c = 36;
      {6'd9, 6'd36} : c = 37;
      {6'd9, 6'd37} : c = 38;
      {6'd9, 6'd38} : c = 39;
      {6'd9, 6'd39} : c = 40;
      {6'd9, 6'd40} : c = 41;
      {6'd9, 6'd41} : c = 42;
      {6'd9, 6'd42} : c = 43;
      {6'd9, 6'd43} : c = 44;
      {6'd9, 6'd44} : c = 45;
      {6'd9, 6'd45} : c = 46;
      {6'd9, 6'd46} : c = 47;
      {6'd9, 6'd47} : c = 48;
      {6'd9, 6'd48} : c = 49;
      {6'd9, 6'd49} : c = 50;
      {6'd9, 6'd50} : c = 51;
      {6'd9, 6'd51} : c = 52;
      {6'd9, 6'd52} : c = 53;
      {6'd9, 6'd53} : c = 54;
      {6'd9, 6'd54} : c = 55;
      {6'd9, 6'd55} : c = 56;
      {6'd9, 6'd56} : c = 57;
      {6'd9, 6'd57} : c = 58;
      {6'd9, 6'd58} : c = 59;
      {6'd9, 6'd59} : c = 60;
      {6'd9, 6'd60} : c = 61;
      {6'd9, 6'd61} : c = 62;
      {6'd9, 6'd62} : c = 63;
      {6'd9, 6'd63} : c = 64;
      {6'd10, 6'd10} : c = 14;
      {6'd10, 6'd11} : c = 15;
      {6'd10, 6'd12} : c = 16;
      {6'd10, 6'd13} : c = 16;
      {6'd10, 6'd14} : c = 17;
      {6'd10, 6'd15} : c = 18;
      {6'd10, 6'd16} : c = 19;
      {6'd10, 6'd17} : c = 20;
      {6'd10, 6'd18} : c = 21;
      {6'd10, 6'd19} : c = 21;
      {6'd10, 6'd20} : c = 22;
      {6'd10, 6'd21} : c = 23;
      {6'd10, 6'd22} : c = 24;
      {6'd10, 6'd23} : c = 25;
      {6'd10, 6'd24} : c = 26;
      {6'd10, 6'd25} : c = 27;
      {6'd10, 6'd26} : c = 28;
      {6'd10, 6'd27} : c = 29;
      {6'd10, 6'd28} : c = 30;
      {6'd10, 6'd29} : c = 31;
      {6'd10, 6'd30} : c = 32;
      {6'd10, 6'd31} : c = 33;
      {6'd10, 6'd32} : c = 34;
      {6'd10, 6'd33} : c = 34;
      {6'd10, 6'd34} : c = 35;
      {6'd10, 6'd35} : c = 36;
      {6'd10, 6'd36} : c = 37;
      {6'd10, 6'd37} : c = 38;
      {6'd10, 6'd38} : c = 39;
      {6'd10, 6'd39} : c = 40;
      {6'd10, 6'd40} : c = 41;
      {6'd10, 6'd41} : c = 42;
      {6'd10, 6'd42} : c = 43;
      {6'd10, 6'd43} : c = 44;
      {6'd10, 6'd44} : c = 45;
      {6'd10, 6'd45} : c = 46;
      {6'd10, 6'd46} : c = 47;
      {6'd10, 6'd47} : c = 48;
      {6'd10, 6'd48} : c = 49;
      {6'd10, 6'd49} : c = 50;
      {6'd10, 6'd50} : c = 51;
      {6'd10, 6'd51} : c = 52;
      {6'd10, 6'd52} : c = 53;
      {6'd10, 6'd53} : c = 54;
      {6'd10, 6'd54} : c = 55;
      {6'd10, 6'd55} : c = 56;
      {6'd10, 6'd56} : c = 57;
      {6'd10, 6'd57} : c = 58;
      {6'd10, 6'd58} : c = 59;
      {6'd10, 6'd59} : c = 60;
      {6'd10, 6'd60} : c = 61;
      {6'd10, 6'd61} : c = 62;
      {6'd10, 6'd62} : c = 63;
      {6'd10, 6'd63} : c = 64;
      {6'd11, 6'd11} : c = 16;
      {6'd11, 6'd12} : c = 16;
      {6'd11, 6'd13} : c = 17;
      {6'd11, 6'd14} : c = 18;
      {6'd11, 6'd15} : c = 19;
      {6'd11, 6'd16} : c = 19;
      {6'd11, 6'd17} : c = 20;
      {6'd11, 6'd18} : c = 21;
      {6'd11, 6'd19} : c = 22;
      {6'd11, 6'd20} : c = 23;
      {6'd11, 6'd21} : c = 24;
      {6'd11, 6'd22} : c = 25;
      {6'd11, 6'd23} : c = 25;
      {6'd11, 6'd24} : c = 26;
      {6'd11, 6'd25} : c = 27;
      {6'd11, 6'd26} : c = 28;
      {6'd11, 6'd27} : c = 29;
      {6'd11, 6'd28} : c = 30;
      {6'd11, 6'd29} : c = 31;
      {6'd11, 6'd30} : c = 32;
      {6'd11, 6'd31} : c = 33;
      {6'd11, 6'd32} : c = 34;
      {6'd11, 6'd33} : c = 35;
      {6'd11, 6'd34} : c = 36;
      {6'd11, 6'd35} : c = 37;
      {6'd11, 6'd36} : c = 38;
      {6'd11, 6'd37} : c = 39;
      {6'd11, 6'd38} : c = 40;
      {6'd11, 6'd39} : c = 41;
      {6'd11, 6'd40} : c = 41;
      {6'd11, 6'd41} : c = 42;
      {6'd11, 6'd42} : c = 43;
      {6'd11, 6'd43} : c = 44;
      {6'd11, 6'd44} : c = 45;
      {6'd11, 6'd45} : c = 46;
      {6'd11, 6'd46} : c = 47;
      {6'd11, 6'd47} : c = 48;
      {6'd11, 6'd48} : c = 49;
      {6'd11, 6'd49} : c = 50;
      {6'd11, 6'd50} : c = 51;
      {6'd11, 6'd51} : c = 52;
      {6'd11, 6'd52} : c = 53;
      {6'd11, 6'd53} : c = 54;
      {6'd11, 6'd54} : c = 55;
      {6'd11, 6'd55} : c = 56;
      {6'd11, 6'd56} : c = 57;
      {6'd11, 6'd57} : c = 58;
      {6'd11, 6'd58} : c = 59;
      {6'd11, 6'd59} : c = 60;
      {6'd11, 6'd60} : c = 61;
      {6'd11, 6'd61} : c = 62;
      {6'd11, 6'd62} : c = 63;
      {6'd11, 6'd63} : c = 64;
      {6'd12, 6'd12} : c = 17;
      {6'd12, 6'd13} : c = 18;
      {6'd12, 6'd14} : c = 18;
      {6'd12, 6'd15} : c = 19;
      {6'd12, 6'd16} : c = 20;
      {6'd12, 6'd17} : c = 21;
      {6'd12, 6'd18} : c = 22;
      {6'd12, 6'd19} : c = 22;
      {6'd12, 6'd20} : c = 23;
      {6'd12, 6'd21} : c = 24;
      {6'd12, 6'd22} : c = 25;
      {6'd12, 6'd23} : c = 26;
      {6'd12, 6'd24} : c = 27;
      {6'd12, 6'd25} : c = 28;
      {6'd12, 6'd26} : c = 29;
      {6'd12, 6'd27} : c = 30;
      {6'd12, 6'd28} : c = 30;
      {6'd12, 6'd29} : c = 31;
      {6'd12, 6'd30} : c = 32;
      {6'd12, 6'd31} : c = 33;
      {6'd12, 6'd32} : c = 34;
      {6'd12, 6'd33} : c = 35;
      {6'd12, 6'd34} : c = 36;
      {6'd12, 6'd35} : c = 37;
      {6'd12, 6'd36} : c = 38;
      {6'd12, 6'd37} : c = 39;
      {6'd12, 6'd38} : c = 40;
      {6'd12, 6'd39} : c = 41;
      {6'd12, 6'd40} : c = 42;
      {6'd12, 6'd41} : c = 43;
      {6'd12, 6'd42} : c = 44;
      {6'd12, 6'd43} : c = 45;
      {6'd12, 6'd44} : c = 46;
      {6'd12, 6'd45} : c = 47;
      {6'd12, 6'd46} : c = 48;
      {6'd12, 6'd47} : c = 49;
      {6'd12, 6'd48} : c = 49;
      {6'd12, 6'd49} : c = 50;
      {6'd12, 6'd50} : c = 51;
      {6'd12, 6'd51} : c = 52;
      {6'd12, 6'd52} : c = 53;
      {6'd12, 6'd53} : c = 54;
      {6'd12, 6'd54} : c = 55;
      {6'd12, 6'd55} : c = 56;
      {6'd12, 6'd56} : c = 57;
      {6'd12, 6'd57} : c = 58;
      {6'd12, 6'd58} : c = 59;
      {6'd12, 6'd59} : c = 60;
      {6'd12, 6'd60} : c = 61;
      {6'd12, 6'd61} : c = 62;
      {6'd12, 6'd62} : c = 63;
      {6'd12, 6'd63} : c = 64;
      {6'd13, 6'd13} : c = 18;
      {6'd13, 6'd14} : c = 19;
      {6'd13, 6'd15} : c = 20;
      {6'd13, 6'd16} : c = 21;
      {6'd13, 6'd17} : c = 21;
      {6'd13, 6'd18} : c = 22;
      {6'd13, 6'd19} : c = 23;
      {6'd13, 6'd20} : c = 24;
      {6'd13, 6'd21} : c = 25;
      {6'd13, 6'd22} : c = 26;
      {6'd13, 6'd23} : c = 26;
      {6'd13, 6'd24} : c = 27;
      {6'd13, 6'd25} : c = 28;
      {6'd13, 6'd26} : c = 29;
      {6'd13, 6'd27} : c = 30;
      {6'd13, 6'd28} : c = 31;
      {6'd13, 6'd29} : c = 32;
      {6'd13, 6'd30} : c = 33;
      {6'd13, 6'd31} : c = 34;
      {6'd13, 6'd32} : c = 35;
      {6'd13, 6'd33} : c = 35;
      {6'd13, 6'd34} : c = 36;
      {6'd13, 6'd35} : c = 37;
      {6'd13, 6'd36} : c = 38;
      {6'd13, 6'd37} : c = 39;
      {6'd13, 6'd38} : c = 40;
      {6'd13, 6'd39} : c = 41;
      {6'd13, 6'd40} : c = 42;
      {6'd13, 6'd41} : c = 43;
      {6'd13, 6'd42} : c = 44;
      {6'd13, 6'd43} : c = 45;
      {6'd13, 6'd44} : c = 46;
      {6'd13, 6'd45} : c = 47;
      {6'd13, 6'd46} : c = 48;
      {6'd13, 6'd47} : c = 49;
      {6'd13, 6'd48} : c = 50;
      {6'd13, 6'd49} : c = 51;
      {6'd13, 6'd50} : c = 52;
      {6'd13, 6'd51} : c = 53;
      {6'd13, 6'd52} : c = 54;
      {6'd13, 6'd53} : c = 55;
      {6'd13, 6'd54} : c = 56;
      {6'd13, 6'd55} : c = 57;
      {6'd13, 6'd56} : c = 57;
      {6'd13, 6'd57} : c = 58;
      {6'd13, 6'd58} : c = 59;
      {6'd13, 6'd59} : c = 60;
      {6'd13, 6'd60} : c = 61;
      {6'd13, 6'd61} : c = 62;
      {6'd13, 6'd62} : c = 63;
      {6'd13, 6'd63} : c = 64;
      {6'd14, 6'd14} : c = 20;
      {6'd14, 6'd15} : c = 21;
      {6'd14, 6'd16} : c = 21;
      {6'd14, 6'd17} : c = 22;
      {6'd14, 6'd18} : c = 23;
      {6'd14, 6'd19} : c = 24;
      {6'd14, 6'd20} : c = 24;
      {6'd14, 6'd21} : c = 25;
      {6'd14, 6'd22} : c = 26;
      {6'd14, 6'd23} : c = 27;
      {6'd14, 6'd24} : c = 28;
      {6'd14, 6'd25} : c = 29;
      {6'd14, 6'd26} : c = 30;
      {6'd14, 6'd27} : c = 30;
      {6'd14, 6'd28} : c = 31;
      {6'd14, 6'd29} : c = 32;
      {6'd14, 6'd30} : c = 33;
      {6'd14, 6'd31} : c = 34;
      {6'd14, 6'd32} : c = 35;
      {6'd14, 6'd33} : c = 36;
      {6'd14, 6'd34} : c = 37;
      {6'd14, 6'd35} : c = 38;
      {6'd14, 6'd36} : c = 39;
      {6'd14, 6'd37} : c = 40;
      {6'd14, 6'd38} : c = 40;
      {6'd14, 6'd39} : c = 41;
      {6'd14, 6'd40} : c = 42;
      {6'd14, 6'd41} : c = 43;
      {6'd14, 6'd42} : c = 44;
      {6'd14, 6'd43} : c = 45;
      {6'd14, 6'd44} : c = 46;
      {6'd14, 6'd45} : c = 47;
      {6'd14, 6'd46} : c = 48;
      {6'd14, 6'd47} : c = 49;
      {6'd14, 6'd48} : c = 50;
      {6'd14, 6'd49} : c = 51;
      {6'd14, 6'd50} : c = 52;
      {6'd14, 6'd51} : c = 53;
      {6'd14, 6'd52} : c = 54;
      {6'd14, 6'd53} : c = 55;
      {6'd14, 6'd54} : c = 56;
      {6'd14, 6'd55} : c = 57;
      {6'd14, 6'd56} : c = 58;
      {6'd14, 6'd57} : c = 59;
      {6'd14, 6'd58} : c = 60;
      {6'd14, 6'd59} : c = 61;
      {6'd14, 6'd60} : c = 62;
      {6'd14, 6'd61} : c = 63;
      {6'd14, 6'd62} : c = 64;
      {6'd14, 6'd63} : c = 65;
      {6'd15, 6'd15} : c = 21;
      {6'd15, 6'd16} : c = 22;
      {6'd15, 6'd17} : c = 23;
      {6'd15, 6'd18} : c = 23;
      {6'd15, 6'd19} : c = 24;
      {6'd15, 6'd20} : c = 25;
      {6'd15, 6'd21} : c = 26;
      {6'd15, 6'd22} : c = 27;
      {6'd15, 6'd23} : c = 27;
      {6'd15, 6'd24} : c = 28;
      {6'd15, 6'd25} : c = 29;
      {6'd15, 6'd26} : c = 30;
      {6'd15, 6'd27} : c = 31;
      {6'd15, 6'd28} : c = 32;
      {6'd15, 6'd29} : c = 33;
      {6'd15, 6'd30} : c = 34;
      {6'd15, 6'd31} : c = 34;
      {6'd15, 6'd32} : c = 35;
      {6'd15, 6'd33} : c = 36;
      {6'd15, 6'd34} : c = 37;
      {6'd15, 6'd35} : c = 38;
      {6'd15, 6'd36} : c = 39;
      {6'd15, 6'd37} : c = 40;
      {6'd15, 6'd38} : c = 41;
      {6'd15, 6'd39} : c = 42;
      {6'd15, 6'd40} : c = 43;
      {6'd15, 6'd41} : c = 44;
      {6'd15, 6'd42} : c = 45;
      {6'd15, 6'd43} : c = 46;
      {6'd15, 6'd44} : c = 46;
      {6'd15, 6'd45} : c = 47;
      {6'd15, 6'd46} : c = 48;
      {6'd15, 6'd47} : c = 49;
      {6'd15, 6'd48} : c = 50;
      {6'd15, 6'd49} : c = 51;
      {6'd15, 6'd50} : c = 52;
      {6'd15, 6'd51} : c = 53;
      {6'd15, 6'd52} : c = 54;
      {6'd15, 6'd53} : c = 55;
      {6'd15, 6'd54} : c = 56;
      {6'd15, 6'd55} : c = 57;
      {6'd15, 6'd56} : c = 58;
      {6'd15, 6'd57} : c = 59;
      {6'd15, 6'd58} : c = 60;
      {6'd15, 6'd59} : c = 61;
      {6'd15, 6'd60} : c = 62;
      {6'd15, 6'd61} : c = 63;
      {6'd15, 6'd62} : c = 64;
      {6'd15, 6'd63} : c = 65;
      {6'd16, 6'd16} : c = 23;
      {6'd16, 6'd17} : c = 23;
      {6'd16, 6'd18} : c = 24;
      {6'd16, 6'd19} : c = 25;
      {6'd16, 6'd20} : c = 26;
      {6'd16, 6'd21} : c = 26;
      {6'd16, 6'd22} : c = 27;
      {6'd16, 6'd23} : c = 28;
      {6'd16, 6'd24} : c = 29;
      {6'd16, 6'd25} : c = 30;
      {6'd16, 6'd26} : c = 31;
      {6'd16, 6'd27} : c = 31;
      {6'd16, 6'd28} : c = 32;
      {6'd16, 6'd29} : c = 33;
      {6'd16, 6'd30} : c = 34;
      {6'd16, 6'd31} : c = 35;
      {6'd16, 6'd32} : c = 36;
      {6'd16, 6'd33} : c = 37;
      {6'd16, 6'd34} : c = 38;
      {6'd16, 6'd35} : c = 38;
      {6'd16, 6'd36} : c = 39;
      {6'd16, 6'd37} : c = 40;
      {6'd16, 6'd38} : c = 41;
      {6'd16, 6'd39} : c = 42;
      {6'd16, 6'd40} : c = 43;
      {6'd16, 6'd41} : c = 44;
      {6'd16, 6'd42} : c = 45;
      {6'd16, 6'd43} : c = 46;
      {6'd16, 6'd44} : c = 47;
      {6'd16, 6'd45} : c = 48;
      {6'd16, 6'd46} : c = 49;
      {6'd16, 6'd47} : c = 50;
      {6'd16, 6'd48} : c = 51;
      {6'd16, 6'd49} : c = 52;
      {6'd16, 6'd50} : c = 52;
      {6'd16, 6'd51} : c = 53;
      {6'd16, 6'd52} : c = 54;
      {6'd16, 6'd53} : c = 55;
      {6'd16, 6'd54} : c = 56;
      {6'd16, 6'd55} : c = 57;
      {6'd16, 6'd56} : c = 58;
      {6'd16, 6'd57} : c = 59;
      {6'd16, 6'd58} : c = 60;
      {6'd16, 6'd59} : c = 61;
      {6'd16, 6'd60} : c = 62;
      {6'd16, 6'd61} : c = 63;
      {6'd16, 6'd62} : c = 64;
      {6'd16, 6'd63} : c = 65;
      {6'd17, 6'd17} : c = 24;
      {6'd17, 6'd18} : c = 25;
      {6'd17, 6'd19} : c = 25;
      {6'd17, 6'd20} : c = 26;
      {6'd17, 6'd21} : c = 27;
      {6'd17, 6'd22} : c = 28;
      {6'd17, 6'd23} : c = 29;
      {6'd17, 6'd24} : c = 29;
      {6'd17, 6'd25} : c = 30;
      {6'd17, 6'd26} : c = 31;
      {6'd17, 6'd27} : c = 32;
      {6'd17, 6'd28} : c = 33;
      {6'd17, 6'd29} : c = 34;
      {6'd17, 6'd30} : c = 34;
      {6'd17, 6'd31} : c = 35;
      {6'd17, 6'd32} : c = 36;
      {6'd17, 6'd33} : c = 37;
      {6'd17, 6'd34} : c = 38;
      {6'd17, 6'd35} : c = 39;
      {6'd17, 6'd36} : c = 40;
      {6'd17, 6'd37} : c = 41;
      {6'd17, 6'd38} : c = 42;
      {6'd17, 6'd39} : c = 43;
      {6'd17, 6'd40} : c = 43;
      {6'd17, 6'd41} : c = 44;
      {6'd17, 6'd42} : c = 45;
      {6'd17, 6'd43} : c = 46;
      {6'd17, 6'd44} : c = 47;
      {6'd17, 6'd45} : c = 48;
      {6'd17, 6'd46} : c = 49;
      {6'd17, 6'd47} : c = 50;
      {6'd17, 6'd48} : c = 51;
      {6'd17, 6'd49} : c = 52;
      {6'd17, 6'd50} : c = 53;
      {6'd17, 6'd51} : c = 54;
      {6'd17, 6'd52} : c = 55;
      {6'd17, 6'd53} : c = 56;
      {6'd17, 6'd54} : c = 57;
      {6'd17, 6'd55} : c = 58;
      {6'd17, 6'd56} : c = 59;
      {6'd17, 6'd57} : c = 59;
      {6'd17, 6'd58} : c = 60;
      {6'd17, 6'd59} : c = 61;
      {6'd17, 6'd60} : c = 62;
      {6'd17, 6'd61} : c = 63;
      {6'd17, 6'd62} : c = 64;
      {6'd17, 6'd63} : c = 65;
      {6'd18, 6'd18} : c = 25;
      {6'd18, 6'd19} : c = 26;
      {6'd18, 6'd20} : c = 27;
      {6'd18, 6'd21} : c = 28;
      {6'd18, 6'd22} : c = 28;
      {6'd18, 6'd23} : c = 29;
      {6'd18, 6'd24} : c = 30;
      {6'd18, 6'd25} : c = 31;
      {6'd18, 6'd26} : c = 32;
      {6'd18, 6'd27} : c = 32;
      {6'd18, 6'd28} : c = 33;
      {6'd18, 6'd29} : c = 34;
      {6'd18, 6'd30} : c = 35;
      {6'd18, 6'd31} : c = 36;
      {6'd18, 6'd32} : c = 37;
      {6'd18, 6'd33} : c = 38;
      {6'd18, 6'd34} : c = 38;
      {6'd18, 6'd35} : c = 39;
      {6'd18, 6'd36} : c = 40;
      {6'd18, 6'd37} : c = 41;
      {6'd18, 6'd38} : c = 42;
      {6'd18, 6'd39} : c = 43;
      {6'd18, 6'd40} : c = 44;
      {6'd18, 6'd41} : c = 45;
      {6'd18, 6'd42} : c = 46;
      {6'd18, 6'd43} : c = 47;
      {6'd18, 6'd44} : c = 48;
      {6'd18, 6'd45} : c = 48;
      {6'd18, 6'd46} : c = 49;
      {6'd18, 6'd47} : c = 50;
      {6'd18, 6'd48} : c = 51;
      {6'd18, 6'd49} : c = 52;
      {6'd18, 6'd50} : c = 53;
      {6'd18, 6'd51} : c = 54;
      {6'd18, 6'd52} : c = 55;
      {6'd18, 6'd53} : c = 56;
      {6'd18, 6'd54} : c = 57;
      {6'd18, 6'd55} : c = 58;
      {6'd18, 6'd56} : c = 59;
      {6'd18, 6'd57} : c = 60;
      {6'd18, 6'd58} : c = 61;
      {6'd18, 6'd59} : c = 62;
      {6'd18, 6'd60} : c = 63;
      {6'd18, 6'd61} : c = 64;
      {6'd18, 6'd62} : c = 65;
      {6'd18, 6'd63} : c = 66;
      {6'd19, 6'd19} : c = 27;
      {6'd19, 6'd20} : c = 28;
      {6'd19, 6'd21} : c = 28;
      {6'd19, 6'd22} : c = 29;
      {6'd19, 6'd23} : c = 30;
      {6'd19, 6'd24} : c = 31;
      {6'd19, 6'd25} : c = 31;
      {6'd19, 6'd26} : c = 32;
      {6'd19, 6'd27} : c = 33;
      {6'd19, 6'd28} : c = 34;
      {6'd19, 6'd29} : c = 35;
      {6'd19, 6'd30} : c = 36;
      {6'd19, 6'd31} : c = 36;
      {6'd19, 6'd32} : c = 37;
      {6'd19, 6'd33} : c = 38;
      {6'd19, 6'd34} : c = 39;
      {6'd19, 6'd35} : c = 40;
      {6'd19, 6'd36} : c = 41;
      {6'd19, 6'd37} : c = 42;
      {6'd19, 6'd38} : c = 42;
      {6'd19, 6'd39} : c = 43;
      {6'd19, 6'd40} : c = 44;
      {6'd19, 6'd41} : c = 45;
      {6'd19, 6'd42} : c = 46;
      {6'd19, 6'd43} : c = 47;
      {6'd19, 6'd44} : c = 48;
      {6'd19, 6'd45} : c = 49;
      {6'd19, 6'd46} : c = 50;
      {6'd19, 6'd47} : c = 51;
      {6'd19, 6'd48} : c = 52;
      {6'd19, 6'd49} : c = 53;
      {6'd19, 6'd50} : c = 53;
      {6'd19, 6'd51} : c = 54;
      {6'd19, 6'd52} : c = 55;
      {6'd19, 6'd53} : c = 56;
      {6'd19, 6'd54} : c = 57;
      {6'd19, 6'd55} : c = 58;
      {6'd19, 6'd56} : c = 59;
      {6'd19, 6'd57} : c = 60;
      {6'd19, 6'd58} : c = 61;
      {6'd19, 6'd59} : c = 62;
      {6'd19, 6'd60} : c = 63;
      {6'd19, 6'd61} : c = 64;
      {6'd19, 6'd62} : c = 65;
      {6'd19, 6'd63} : c = 66;
      {6'd20, 6'd20} : c = 28;
      {6'd20, 6'd21} : c = 29;
      {6'd20, 6'd22} : c = 30;
      {6'd20, 6'd23} : c = 30;
      {6'd20, 6'd24} : c = 31;
      {6'd20, 6'd25} : c = 32;
      {6'd20, 6'd26} : c = 33;
      {6'd20, 6'd27} : c = 34;
      {6'd20, 6'd28} : c = 34;
      {6'd20, 6'd29} : c = 35;
      {6'd20, 6'd30} : c = 36;
      {6'd20, 6'd31} : c = 37;
      {6'd20, 6'd32} : c = 38;
      {6'd20, 6'd33} : c = 39;
      {6'd20, 6'd34} : c = 39;
      {6'd20, 6'd35} : c = 40;
      {6'd20, 6'd36} : c = 41;
      {6'd20, 6'd37} : c = 42;
      {6'd20, 6'd38} : c = 43;
      {6'd20, 6'd39} : c = 44;
      {6'd20, 6'd40} : c = 45;
      {6'd20, 6'd41} : c = 46;
      {6'd20, 6'd42} : c = 47;
      {6'd20, 6'd43} : c = 47;
      {6'd20, 6'd44} : c = 48;
      {6'd20, 6'd45} : c = 49;
      {6'd20, 6'd46} : c = 50;
      {6'd20, 6'd47} : c = 51;
      {6'd20, 6'd48} : c = 52;
      {6'd20, 6'd49} : c = 53;
      {6'd20, 6'd50} : c = 54;
      {6'd20, 6'd51} : c = 55;
      {6'd20, 6'd52} : c = 56;
      {6'd20, 6'd53} : c = 57;
      {6'd20, 6'd54} : c = 58;
      {6'd20, 6'd55} : c = 59;
      {6'd20, 6'd56} : c = 59;
      {6'd20, 6'd57} : c = 60;
      {6'd20, 6'd58} : c = 61;
      {6'd20, 6'd59} : c = 62;
      {6'd20, 6'd60} : c = 63;
      {6'd20, 6'd61} : c = 64;
      {6'd20, 6'd62} : c = 65;
      {6'd20, 6'd63} : c = 66;
      {6'd21, 6'd21} : c = 30;
      {6'd21, 6'd22} : c = 30;
      {6'd21, 6'd23} : c = 31;
      {6'd21, 6'd24} : c = 32;
      {6'd21, 6'd25} : c = 33;
      {6'd21, 6'd26} : c = 33;
      {6'd21, 6'd27} : c = 34;
      {6'd21, 6'd28} : c = 35;
      {6'd21, 6'd29} : c = 36;
      {6'd21, 6'd30} : c = 37;
      {6'd21, 6'd31} : c = 37;
      {6'd21, 6'd32} : c = 38;
      {6'd21, 6'd33} : c = 39;
      {6'd21, 6'd34} : c = 40;
      {6'd21, 6'd35} : c = 41;
      {6'd21, 6'd36} : c = 42;
      {6'd21, 6'd37} : c = 43;
      {6'd21, 6'd38} : c = 43;
      {6'd21, 6'd39} : c = 44;
      {6'd21, 6'd40} : c = 45;
      {6'd21, 6'd41} : c = 46;
      {6'd21, 6'd42} : c = 47;
      {6'd21, 6'd43} : c = 48;
      {6'd21, 6'd44} : c = 49;
      {6'd21, 6'd45} : c = 50;
      {6'd21, 6'd46} : c = 51;
      {6'd21, 6'd47} : c = 51;
      {6'd21, 6'd48} : c = 52;
      {6'd21, 6'd49} : c = 53;
      {6'd21, 6'd50} : c = 54;
      {6'd21, 6'd51} : c = 55;
      {6'd21, 6'd52} : c = 56;
      {6'd21, 6'd53} : c = 57;
      {6'd21, 6'd54} : c = 58;
      {6'd21, 6'd55} : c = 59;
      {6'd21, 6'd56} : c = 60;
      {6'd21, 6'd57} : c = 61;
      {6'd21, 6'd58} : c = 62;
      {6'd21, 6'd59} : c = 63;
      {6'd21, 6'd60} : c = 64;
      {6'd21, 6'd61} : c = 65;
      {6'd21, 6'd62} : c = 65;
      {6'd21, 6'd63} : c = 66;
      {6'd22, 6'd22} : c = 31;
      {6'd22, 6'd23} : c = 32;
      {6'd22, 6'd24} : c = 33;
      {6'd22, 6'd25} : c = 33;
      {6'd22, 6'd26} : c = 34;
      {6'd22, 6'd27} : c = 35;
      {6'd22, 6'd28} : c = 36;
      {6'd22, 6'd29} : c = 36;
      {6'd22, 6'd30} : c = 37;
      {6'd22, 6'd31} : c = 38;
      {6'd22, 6'd32} : c = 39;
      {6'd22, 6'd33} : c = 40;
      {6'd22, 6'd34} : c = 40;
      {6'd22, 6'd35} : c = 41;
      {6'd22, 6'd36} : c = 42;
      {6'd22, 6'd37} : c = 43;
      {6'd22, 6'd38} : c = 44;
      {6'd22, 6'd39} : c = 45;
      {6'd22, 6'd40} : c = 46;
      {6'd22, 6'd41} : c = 47;
      {6'd22, 6'd42} : c = 47;
      {6'd22, 6'd43} : c = 48;
      {6'd22, 6'd44} : c = 49;
      {6'd22, 6'd45} : c = 50;
      {6'd22, 6'd46} : c = 51;
      {6'd22, 6'd47} : c = 52;
      {6'd22, 6'd48} : c = 53;
      {6'd22, 6'd49} : c = 54;
      {6'd22, 6'd50} : c = 55;
      {6'd22, 6'd51} : c = 56;
      {6'd22, 6'd52} : c = 56;
      {6'd22, 6'd53} : c = 57;
      {6'd22, 6'd54} : c = 58;
      {6'd22, 6'd55} : c = 59;
      {6'd22, 6'd56} : c = 60;
      {6'd22, 6'd57} : c = 61;
      {6'd22, 6'd58} : c = 62;
      {6'd22, 6'd59} : c = 63;
      {6'd22, 6'd60} : c = 64;
      {6'd22, 6'd61} : c = 65;
      {6'd22, 6'd62} : c = 66;
      {6'd22, 6'd63} : c = 67;
      {6'd23, 6'd23} : c = 33;
      {6'd23, 6'd24} : c = 33;
      {6'd23, 6'd25} : c = 34;
      {6'd23, 6'd26} : c = 35;
      {6'd23, 6'd27} : c = 35;
      {6'd23, 6'd28} : c = 36;
      {6'd23, 6'd29} : c = 37;
      {6'd23, 6'd30} : c = 38;
      {6'd23, 6'd31} : c = 39;
      {6'd23, 6'd32} : c = 39;
      {6'd23, 6'd33} : c = 40;
      {6'd23, 6'd34} : c = 41;
      {6'd23, 6'd35} : c = 42;
      {6'd23, 6'd36} : c = 43;
      {6'd23, 6'd37} : c = 44;
      {6'd23, 6'd38} : c = 44;
      {6'd23, 6'd39} : c = 45;
      {6'd23, 6'd40} : c = 46;
      {6'd23, 6'd41} : c = 47;
      {6'd23, 6'd42} : c = 48;
      {6'd23, 6'd43} : c = 49;
      {6'd23, 6'd44} : c = 50;
      {6'd23, 6'd45} : c = 51;
      {6'd23, 6'd46} : c = 51;
      {6'd23, 6'd47} : c = 52;
      {6'd23, 6'd48} : c = 53;
      {6'd23, 6'd49} : c = 54;
      {6'd23, 6'd50} : c = 55;
      {6'd23, 6'd51} : c = 56;
      {6'd23, 6'd52} : c = 57;
      {6'd23, 6'd53} : c = 58;
      {6'd23, 6'd54} : c = 59;
      {6'd23, 6'd55} : c = 60;
      {6'd23, 6'd56} : c = 61;
      {6'd23, 6'd57} : c = 61;
      {6'd23, 6'd58} : c = 62;
      {6'd23, 6'd59} : c = 63;
      {6'd23, 6'd60} : c = 64;
      {6'd23, 6'd61} : c = 65;
      {6'd23, 6'd62} : c = 66;
      {6'd23, 6'd63} : c = 67;
      {6'd24, 6'd24} : c = 34;
      {6'd24, 6'd25} : c = 35;
      {6'd24, 6'd26} : c = 35;
      {6'd24, 6'd27} : c = 36;
      {6'd24, 6'd28} : c = 37;
      {6'd24, 6'd29} : c = 38;
      {6'd24, 6'd30} : c = 38;
      {6'd24, 6'd31} : c = 39;
      {6'd24, 6'd32} : c = 40;
      {6'd24, 6'd33} : c = 41;
      {6'd24, 6'd34} : c = 42;
      {6'd24, 6'd35} : c = 42;
      {6'd24, 6'd36} : c = 43;
      {6'd24, 6'd37} : c = 44;
      {6'd24, 6'd38} : c = 45;
      {6'd24, 6'd39} : c = 46;
      {6'd24, 6'd40} : c = 47;
      {6'd24, 6'd41} : c = 48;
      {6'd24, 6'd42} : c = 48;
      {6'd24, 6'd43} : c = 49;
      {6'd24, 6'd44} : c = 50;
      {6'd24, 6'd45} : c = 51;
      {6'd24, 6'd46} : c = 52;
      {6'd24, 6'd47} : c = 53;
      {6'd24, 6'd48} : c = 54;
      {6'd24, 6'd49} : c = 55;
      {6'd24, 6'd50} : c = 55;
      {6'd24, 6'd51} : c = 56;
      {6'd24, 6'd52} : c = 57;
      {6'd24, 6'd53} : c = 58;
      {6'd24, 6'd54} : c = 59;
      {6'd24, 6'd55} : c = 60;
      {6'd24, 6'd56} : c = 61;
      {6'd24, 6'd57} : c = 62;
      {6'd24, 6'd58} : c = 63;
      {6'd24, 6'd59} : c = 64;
      {6'd24, 6'd60} : c = 65;
      {6'd24, 6'd61} : c = 66;
      {6'd24, 6'd62} : c = 66;
      {6'd24, 6'd63} : c = 67;
      {6'd25, 6'd25} : c = 35;
      {6'd25, 6'd26} : c = 36;
      {6'd25, 6'd27} : c = 37;
      {6'd25, 6'd28} : c = 38;
      {6'd25, 6'd29} : c = 38;
      {6'd25, 6'd30} : c = 39;
      {6'd25, 6'd31} : c = 40;
      {6'd25, 6'd32} : c = 41;
      {6'd25, 6'd33} : c = 41;
      {6'd25, 6'd34} : c = 42;
      {6'd25, 6'd35} : c = 43;
      {6'd25, 6'd36} : c = 44;
      {6'd25, 6'd37} : c = 45;
      {6'd25, 6'd38} : c = 45;
      {6'd25, 6'd39} : c = 46;
      {6'd25, 6'd40} : c = 47;
      {6'd25, 6'd41} : c = 48;
      {6'd25, 6'd42} : c = 49;
      {6'd25, 6'd43} : c = 50;
      {6'd25, 6'd44} : c = 51;
      {6'd25, 6'd45} : c = 51;
      {6'd25, 6'd46} : c = 52;
      {6'd25, 6'd47} : c = 53;
      {6'd25, 6'd48} : c = 54;
      {6'd25, 6'd49} : c = 55;
      {6'd25, 6'd50} : c = 56;
      {6'd25, 6'd51} : c = 57;
      {6'd25, 6'd52} : c = 58;
      {6'd25, 6'd53} : c = 59;
      {6'd25, 6'd54} : c = 60;
      {6'd25, 6'd55} : c = 60;
      {6'd25, 6'd56} : c = 61;
      {6'd25, 6'd57} : c = 62;
      {6'd25, 6'd58} : c = 63;
      {6'd25, 6'd59} : c = 64;
      {6'd25, 6'd60} : c = 65;
      {6'd25, 6'd61} : c = 66;
      {6'd25, 6'd62} : c = 67;
      {6'd25, 6'd63} : c = 68;
      {6'd26, 6'd26} : c = 37;
      {6'd26, 6'd27} : c = 37;
      {6'd26, 6'd28} : c = 38;
      {6'd26, 6'd29} : c = 39;
      {6'd26, 6'd30} : c = 40;
      {6'd26, 6'd31} : c = 40;
      {6'd26, 6'd32} : c = 41;
      {6'd26, 6'd33} : c = 42;
      {6'd26, 6'd34} : c = 43;
      {6'd26, 6'd35} : c = 44;
      {6'd26, 6'd36} : c = 44;
      {6'd26, 6'd37} : c = 45;
      {6'd26, 6'd38} : c = 46;
      {6'd26, 6'd39} : c = 47;
      {6'd26, 6'd40} : c = 48;
      {6'd26, 6'd41} : c = 49;
      {6'd26, 6'd42} : c = 49;
      {6'd26, 6'd43} : c = 50;
      {6'd26, 6'd44} : c = 51;
      {6'd26, 6'd45} : c = 52;
      {6'd26, 6'd46} : c = 53;
      {6'd26, 6'd47} : c = 54;
      {6'd26, 6'd48} : c = 55;
      {6'd26, 6'd49} : c = 55;
      {6'd26, 6'd50} : c = 56;
      {6'd26, 6'd51} : c = 57;
      {6'd26, 6'd52} : c = 58;
      {6'd26, 6'd53} : c = 59;
      {6'd26, 6'd54} : c = 60;
      {6'd26, 6'd55} : c = 61;
      {6'd26, 6'd56} : c = 62;
      {6'd26, 6'd57} : c = 63;
      {6'd26, 6'd58} : c = 64;
      {6'd26, 6'd59} : c = 64;
      {6'd26, 6'd60} : c = 65;
      {6'd26, 6'd61} : c = 66;
      {6'd26, 6'd62} : c = 67;
      {6'd26, 6'd63} : c = 68;
      {6'd27, 6'd27} : c = 38;
      {6'd27, 6'd28} : c = 39;
      {6'd27, 6'd29} : c = 40;
      {6'd27, 6'd30} : c = 40;
      {6'd27, 6'd31} : c = 41;
      {6'd27, 6'd32} : c = 42;
      {6'd27, 6'd33} : c = 43;
      {6'd27, 6'd34} : c = 43;
      {6'd27, 6'd35} : c = 44;
      {6'd27, 6'd36} : c = 45;
      {6'd27, 6'd37} : c = 46;
      {6'd27, 6'd38} : c = 47;
      {6'd27, 6'd39} : c = 47;
      {6'd27, 6'd40} : c = 48;
      {6'd27, 6'd41} : c = 49;
      {6'd27, 6'd42} : c = 50;
      {6'd27, 6'd43} : c = 51;
      {6'd27, 6'd44} : c = 52;
      {6'd27, 6'd45} : c = 52;
      {6'd27, 6'd46} : c = 53;
      {6'd27, 6'd47} : c = 54;
      {6'd27, 6'd48} : c = 55;
      {6'd27, 6'd49} : c = 56;
      {6'd27, 6'd50} : c = 57;
      {6'd27, 6'd51} : c = 58;
      {6'd27, 6'd52} : c = 59;
      {6'd27, 6'd53} : c = 59;
      {6'd27, 6'd54} : c = 60;
      {6'd27, 6'd55} : c = 61;
      {6'd27, 6'd56} : c = 62;
      {6'd27, 6'd57} : c = 63;
      {6'd27, 6'd58} : c = 64;
      {6'd27, 6'd59} : c = 65;
      {6'd27, 6'd60} : c = 66;
      {6'd27, 6'd61} : c = 67;
      {6'd27, 6'd62} : c = 68;
      {6'd27, 6'd63} : c = 69;
      {6'd28, 6'd28} : c = 40;
      {6'd28, 6'd29} : c = 40;
      {6'd28, 6'd30} : c = 41;
      {6'd28, 6'd31} : c = 42;
      {6'd28, 6'd32} : c = 43;
      {6'd28, 6'd33} : c = 43;
      {6'd28, 6'd34} : c = 44;
      {6'd28, 6'd35} : c = 45;
      {6'd28, 6'd36} : c = 46;
      {6'd28, 6'd37} : c = 46;
      {6'd28, 6'd38} : c = 47;
      {6'd28, 6'd39} : c = 48;
      {6'd28, 6'd40} : c = 49;
      {6'd28, 6'd41} : c = 50;
      {6'd28, 6'd42} : c = 50;
      {6'd28, 6'd43} : c = 51;
      {6'd28, 6'd44} : c = 52;
      {6'd28, 6'd45} : c = 53;
      {6'd28, 6'd46} : c = 54;
      {6'd28, 6'd47} : c = 55;
      {6'd28, 6'd48} : c = 56;
      {6'd28, 6'd49} : c = 56;
      {6'd28, 6'd50} : c = 57;
      {6'd28, 6'd51} : c = 58;
      {6'd28, 6'd52} : c = 59;
      {6'd28, 6'd53} : c = 60;
      {6'd28, 6'd54} : c = 61;
      {6'd28, 6'd55} : c = 62;
      {6'd28, 6'd56} : c = 63;
      {6'd28, 6'd57} : c = 64;
      {6'd28, 6'd58} : c = 64;
      {6'd28, 6'd59} : c = 65;
      {6'd28, 6'd60} : c = 66;
      {6'd28, 6'd61} : c = 67;
      {6'd28, 6'd62} : c = 68;
      {6'd28, 6'd63} : c = 69;
      {6'd29, 6'd29} : c = 41;
      {6'd29, 6'd30} : c = 42;
      {6'd29, 6'd31} : c = 42;
      {6'd29, 6'd32} : c = 43;
      {6'd29, 6'd33} : c = 44;
      {6'd29, 6'd34} : c = 45;
      {6'd29, 6'd35} : c = 45;
      {6'd29, 6'd36} : c = 46;
      {6'd29, 6'd37} : c = 47;
      {6'd29, 6'd38} : c = 48;
      {6'd29, 6'd39} : c = 49;
      {6'd29, 6'd40} : c = 49;
      {6'd29, 6'd41} : c = 50;
      {6'd29, 6'd42} : c = 51;
      {6'd29, 6'd43} : c = 52;
      {6'd29, 6'd44} : c = 53;
      {6'd29, 6'd45} : c = 54;
      {6'd29, 6'd46} : c = 54;
      {6'd29, 6'd47} : c = 55;
      {6'd29, 6'd48} : c = 56;
      {6'd29, 6'd49} : c = 57;
      {6'd29, 6'd50} : c = 58;
      {6'd29, 6'd51} : c = 59;
      {6'd29, 6'd52} : c = 60;
      {6'd29, 6'd53} : c = 60;
      {6'd29, 6'd54} : c = 61;
      {6'd29, 6'd55} : c = 62;
      {6'd29, 6'd56} : c = 63;
      {6'd29, 6'd57} : c = 64;
      {6'd29, 6'd58} : c = 65;
      {6'd29, 6'd59} : c = 66;
      {6'd29, 6'd60} : c = 67;
      {6'd29, 6'd61} : c = 68;
      {6'd29, 6'd62} : c = 68;
      {6'd29, 6'd63} : c = 69;
      {6'd30, 6'd30} : c = 42;
      {6'd30, 6'd31} : c = 43;
      {6'd30, 6'd32} : c = 44;
      {6'd30, 6'd33} : c = 45;
      {6'd30, 6'd34} : c = 45;
      {6'd30, 6'd35} : c = 46;
      {6'd30, 6'd36} : c = 47;
      {6'd30, 6'd37} : c = 48;
      {6'd30, 6'd38} : c = 48;
      {6'd30, 6'd39} : c = 49;
      {6'd30, 6'd40} : c = 50;
      {6'd30, 6'd41} : c = 51;
      {6'd30, 6'd42} : c = 52;
      {6'd30, 6'd43} : c = 52;
      {6'd30, 6'd44} : c = 53;
      {6'd30, 6'd45} : c = 54;
      {6'd30, 6'd46} : c = 55;
      {6'd30, 6'd47} : c = 56;
      {6'd30, 6'd48} : c = 57;
      {6'd30, 6'd49} : c = 57;
      {6'd30, 6'd50} : c = 58;
      {6'd30, 6'd51} : c = 59;
      {6'd30, 6'd52} : c = 60;
      {6'd30, 6'd53} : c = 61;
      {6'd30, 6'd54} : c = 62;
      {6'd30, 6'd55} : c = 63;
      {6'd30, 6'd56} : c = 64;
      {6'd30, 6'd57} : c = 64;
      {6'd30, 6'd58} : c = 65;
      {6'd30, 6'd59} : c = 66;
      {6'd30, 6'd60} : c = 67;
      {6'd30, 6'd61} : c = 68;
      {6'd30, 6'd62} : c = 69;
      {6'd30, 6'd63} : c = 70;
      {6'd31, 6'd31} : c = 44;
      {6'd31, 6'd32} : c = 45;
      {6'd31, 6'd33} : c = 45;
      {6'd31, 6'd34} : c = 46;
      {6'd31, 6'd35} : c = 47;
      {6'd31, 6'd36} : c = 48;
      {6'd31, 6'd37} : c = 48;
      {6'd31, 6'd38} : c = 49;
      {6'd31, 6'd39} : c = 50;
      {6'd31, 6'd40} : c = 51;
      {6'd31, 6'd41} : c = 51;
      {6'd31, 6'd42} : c = 52;
      {6'd31, 6'd43} : c = 53;
      {6'd31, 6'd44} : c = 54;
      {6'd31, 6'd45} : c = 55;
      {6'd31, 6'd46} : c = 55;
      {6'd31, 6'd47} : c = 56;
      {6'd31, 6'd48} : c = 57;
      {6'd31, 6'd49} : c = 58;
      {6'd31, 6'd50} : c = 59;
      {6'd31, 6'd51} : c = 60;
      {6'd31, 6'd52} : c = 61;
      {6'd31, 6'd53} : c = 61;
      {6'd31, 6'd54} : c = 62;
      {6'd31, 6'd55} : c = 63;
      {6'd31, 6'd56} : c = 64;
      {6'd31, 6'd57} : c = 65;
      {6'd31, 6'd58} : c = 66;
      {6'd31, 6'd59} : c = 67;
      {6'd31, 6'd60} : c = 68;
      {6'd31, 6'd61} : c = 68;
      {6'd31, 6'd62} : c = 69;
      {6'd31, 6'd63} : c = 70;
      {6'd32, 6'd32} : c = 45;
      {6'd32, 6'd33} : c = 46;
      {6'd32, 6'd34} : c = 47;
      {6'd32, 6'd35} : c = 47;
      {6'd32, 6'd36} : c = 48;
      {6'd32, 6'd37} : c = 49;
      {6'd32, 6'd38} : c = 50;
      {6'd32, 6'd39} : c = 50;
      {6'd32, 6'd40} : c = 51;
      {6'd32, 6'd41} : c = 52;
      {6'd32, 6'd42} : c = 53;
      {6'd32, 6'd43} : c = 54;
      {6'd32, 6'd44} : c = 54;
      {6'd32, 6'd45} : c = 55;
      {6'd32, 6'd46} : c = 56;
      {6'd32, 6'd47} : c = 57;
      {6'd32, 6'd48} : c = 58;
      {6'd32, 6'd49} : c = 59;
      {6'd32, 6'd50} : c = 59;
      {6'd32, 6'd51} : c = 60;
      {6'd32, 6'd52} : c = 61;
      {6'd32, 6'd53} : c = 62;
      {6'd32, 6'd54} : c = 63;
      {6'd32, 6'd55} : c = 64;
      {6'd32, 6'd56} : c = 64;
      {6'd32, 6'd57} : c = 65;
      {6'd32, 6'd58} : c = 66;
      {6'd32, 6'd59} : c = 67;
      {6'd32, 6'd60} : c = 68;
      {6'd32, 6'd61} : c = 69;
      {6'd32, 6'd62} : c = 70;
      {6'd32, 6'd63} : c = 71;
      {6'd33, 6'd33} : c = 47;
      {6'd33, 6'd34} : c = 47;
      {6'd33, 6'd35} : c = 48;
      {6'd33, 6'd36} : c = 49;
      {6'd33, 6'd37} : c = 50;
      {6'd33, 6'd38} : c = 50;
      {6'd33, 6'd39} : c = 51;
      {6'd33, 6'd40} : c = 52;
      {6'd33, 6'd41} : c = 53;
      {6'd33, 6'd42} : c = 53;
      {6'd33, 6'd43} : c = 54;
      {6'd33, 6'd44} : c = 55;
      {6'd33, 6'd45} : c = 56;
      {6'd33, 6'd46} : c = 57;
      {6'd33, 6'd47} : c = 57;
      {6'd33, 6'd48} : c = 58;
      {6'd33, 6'd49} : c = 59;
      {6'd33, 6'd50} : c = 60;
      {6'd33, 6'd51} : c = 61;
      {6'd33, 6'd52} : c = 62;
      {6'd33, 6'd53} : c = 62;
      {6'd33, 6'd54} : c = 63;
      {6'd33, 6'd55} : c = 64;
      {6'd33, 6'd56} : c = 65;
      {6'd33, 6'd57} : c = 66;
      {6'd33, 6'd58} : c = 67;
      {6'd33, 6'd59} : c = 68;
      {6'd33, 6'd60} : c = 68;
      {6'd33, 6'd61} : c = 69;
      {6'd33, 6'd62} : c = 70;
      {6'd33, 6'd63} : c = 71;
      {6'd34, 6'd34} : c = 48;
      {6'd34, 6'd35} : c = 49;
      {6'd34, 6'd36} : c = 50;
      {6'd34, 6'd37} : c = 50;
      {6'd34, 6'd38} : c = 51;
      {6'd34, 6'd39} : c = 52;
      {6'd34, 6'd40} : c = 52;
      {6'd34, 6'd41} : c = 53;
      {6'd34, 6'd42} : c = 54;
      {6'd34, 6'd43} : c = 55;
      {6'd34, 6'd44} : c = 56;
      {6'd34, 6'd45} : c = 56;
      {6'd34, 6'd46} : c = 57;
      {6'd34, 6'd47} : c = 58;
      {6'd34, 6'd48} : c = 59;
      {6'd34, 6'd49} : c = 60;
      {6'd34, 6'd50} : c = 60;
      {6'd34, 6'd51} : c = 61;
      {6'd34, 6'd52} : c = 62;
      {6'd34, 6'd53} : c = 63;
      {6'd34, 6'd54} : c = 64;
      {6'd34, 6'd55} : c = 65;
      {6'd34, 6'd56} : c = 66;
      {6'd34, 6'd57} : c = 66;
      {6'd34, 6'd58} : c = 67;
      {6'd34, 6'd59} : c = 68;
      {6'd34, 6'd60} : c = 69;
      {6'd34, 6'd61} : c = 70;
      {6'd34, 6'd62} : c = 71;
      {6'd34, 6'd63} : c = 72;
      {6'd35, 6'd35} : c = 49;
      {6'd35, 6'd36} : c = 50;
      {6'd35, 6'd37} : c = 51;
      {6'd35, 6'd38} : c = 52;
      {6'd35, 6'd39} : c = 52;
      {6'd35, 6'd40} : c = 53;
      {6'd35, 6'd41} : c = 54;
      {6'd35, 6'd42} : c = 55;
      {6'd35, 6'd43} : c = 55;
      {6'd35, 6'd44} : c = 56;
      {6'd35, 6'd45} : c = 57;
      {6'd35, 6'd46} : c = 58;
      {6'd35, 6'd47} : c = 59;
      {6'd35, 6'd48} : c = 59;
      {6'd35, 6'd49} : c = 60;
      {6'd35, 6'd50} : c = 61;
      {6'd35, 6'd51} : c = 62;
      {6'd35, 6'd52} : c = 63;
      {6'd35, 6'd53} : c = 64;
      {6'd35, 6'd54} : c = 64;
      {6'd35, 6'd55} : c = 65;
      {6'd35, 6'd56} : c = 66;
      {6'd35, 6'd57} : c = 67;
      {6'd35, 6'd58} : c = 68;
      {6'd35, 6'd59} : c = 69;
      {6'd35, 6'd60} : c = 69;
      {6'd35, 6'd61} : c = 70;
      {6'd35, 6'd62} : c = 71;
      {6'd35, 6'd63} : c = 72;
      {6'd36, 6'd36} : c = 51;
      {6'd36, 6'd37} : c = 52;
      {6'd36, 6'd38} : c = 52;
      {6'd36, 6'd39} : c = 53;
      {6'd36, 6'd40} : c = 54;
      {6'd36, 6'd41} : c = 55;
      {6'd36, 6'd42} : c = 55;
      {6'd36, 6'd43} : c = 56;
      {6'd36, 6'd44} : c = 57;
      {6'd36, 6'd45} : c = 58;
      {6'd36, 6'd46} : c = 58;
      {6'd36, 6'd47} : c = 59;
      {6'd36, 6'd48} : c = 60;
      {6'd36, 6'd49} : c = 61;
      {6'd36, 6'd50} : c = 62;
      {6'd36, 6'd51} : c = 62;
      {6'd36, 6'd52} : c = 63;
      {6'd36, 6'd53} : c = 64;
      {6'd36, 6'd54} : c = 65;
      {6'd36, 6'd55} : c = 66;
      {6'd36, 6'd56} : c = 67;
      {6'd36, 6'd57} : c = 67;
      {6'd36, 6'd58} : c = 68;
      {6'd36, 6'd59} : c = 69;
      {6'd36, 6'd60} : c = 70;
      {6'd36, 6'd61} : c = 71;
      {6'd36, 6'd62} : c = 72;
      {6'd36, 6'd63} : c = 73;
      {6'd37, 6'd37} : c = 52;
      {6'd37, 6'd38} : c = 53;
      {6'd37, 6'd39} : c = 54;
      {6'd37, 6'd40} : c = 54;
      {6'd37, 6'd41} : c = 55;
      {6'd37, 6'd42} : c = 56;
      {6'd37, 6'd43} : c = 57;
      {6'd37, 6'd44} : c = 57;
      {6'd37, 6'd45} : c = 58;
      {6'd37, 6'd46} : c = 59;
      {6'd37, 6'd47} : c = 60;
      {6'd37, 6'd48} : c = 61;
      {6'd37, 6'd49} : c = 61;
      {6'd37, 6'd50} : c = 62;
      {6'd37, 6'd51} : c = 63;
      {6'd37, 6'd52} : c = 64;
      {6'd37, 6'd53} : c = 65;
      {6'd37, 6'd54} : c = 65;
      {6'd37, 6'd55} : c = 66;
      {6'd37, 6'd56} : c = 67;
      {6'd37, 6'd57} : c = 68;
      {6'd37, 6'd58} : c = 69;
      {6'd37, 6'd59} : c = 70;
      {6'd37, 6'd60} : c = 70;
      {6'd37, 6'd61} : c = 71;
      {6'd37, 6'd62} : c = 72;
      {6'd37, 6'd63} : c = 73;
      {6'd38, 6'd38} : c = 54;
      {6'd38, 6'd39} : c = 54;
      {6'd38, 6'd40} : c = 55;
      {6'd38, 6'd41} : c = 56;
      {6'd38, 6'd42} : c = 57;
      {6'd38, 6'd43} : c = 57;
      {6'd38, 6'd44} : c = 58;
      {6'd38, 6'd45} : c = 59;
      {6'd38, 6'd46} : c = 60;
      {6'd38, 6'd47} : c = 60;
      {6'd38, 6'd48} : c = 61;
      {6'd38, 6'd49} : c = 62;
      {6'd38, 6'd50} : c = 63;
      {6'd38, 6'd51} : c = 64;
      {6'd38, 6'd52} : c = 64;
      {6'd38, 6'd53} : c = 65;
      {6'd38, 6'd54} : c = 66;
      {6'd38, 6'd55} : c = 67;
      {6'd38, 6'd56} : c = 68;
      {6'd38, 6'd57} : c = 69;
      {6'd38, 6'd58} : c = 69;
      {6'd38, 6'd59} : c = 70;
      {6'd38, 6'd60} : c = 71;
      {6'd38, 6'd61} : c = 72;
      {6'd38, 6'd62} : c = 73;
      {6'd38, 6'd63} : c = 74;
      {6'd39, 6'd39} : c = 55;
      {6'd39, 6'd40} : c = 56;
      {6'd39, 6'd41} : c = 57;
      {6'd39, 6'd42} : c = 57;
      {6'd39, 6'd43} : c = 58;
      {6'd39, 6'd44} : c = 59;
      {6'd39, 6'd45} : c = 60;
      {6'd39, 6'd46} : c = 60;
      {6'd39, 6'd47} : c = 61;
      {6'd39, 6'd48} : c = 62;
      {6'd39, 6'd49} : c = 63;
      {6'd39, 6'd50} : c = 63;
      {6'd39, 6'd51} : c = 64;
      {6'd39, 6'd52} : c = 65;
      {6'd39, 6'd53} : c = 66;
      {6'd39, 6'd54} : c = 67;
      {6'd39, 6'd55} : c = 67;
      {6'd39, 6'd56} : c = 68;
      {6'd39, 6'd57} : c = 69;
      {6'd39, 6'd58} : c = 70;
      {6'd39, 6'd59} : c = 71;
      {6'd39, 6'd60} : c = 72;
      {6'd39, 6'd61} : c = 72;
      {6'd39, 6'd62} : c = 73;
      {6'd39, 6'd63} : c = 74;
      {6'd40, 6'd40} : c = 57;
      {6'd40, 6'd41} : c = 57;
      {6'd40, 6'd42} : c = 58;
      {6'd40, 6'd43} : c = 59;
      {6'd40, 6'd44} : c = 59;
      {6'd40, 6'd45} : c = 60;
      {6'd40, 6'd46} : c = 61;
      {6'd40, 6'd47} : c = 62;
      {6'd40, 6'd48} : c = 62;
      {6'd40, 6'd49} : c = 63;
      {6'd40, 6'd50} : c = 64;
      {6'd40, 6'd51} : c = 65;
      {6'd40, 6'd52} : c = 66;
      {6'd40, 6'd53} : c = 66;
      {6'd40, 6'd54} : c = 67;
      {6'd40, 6'd55} : c = 68;
      {6'd40, 6'd56} : c = 69;
      {6'd40, 6'd57} : c = 70;
      {6'd40, 6'd58} : c = 70;
      {6'd40, 6'd59} : c = 71;
      {6'd40, 6'd60} : c = 72;
      {6'd40, 6'd61} : c = 73;
      {6'd40, 6'd62} : c = 74;
      {6'd40, 6'd63} : c = 75;
      {6'd41, 6'd41} : c = 58;
      {6'd41, 6'd42} : c = 59;
      {6'd41, 6'd43} : c = 59;
      {6'd41, 6'd44} : c = 60;
      {6'd41, 6'd45} : c = 61;
      {6'd41, 6'd46} : c = 62;
      {6'd41, 6'd47} : c = 62;
      {6'd41, 6'd48} : c = 63;
      {6'd41, 6'd49} : c = 64;
      {6'd41, 6'd50} : c = 65;
      {6'd41, 6'd51} : c = 65;
      {6'd41, 6'd52} : c = 66;
      {6'd41, 6'd53} : c = 67;
      {6'd41, 6'd54} : c = 68;
      {6'd41, 6'd55} : c = 69;
      {6'd41, 6'd56} : c = 69;
      {6'd41, 6'd57} : c = 70;
      {6'd41, 6'd58} : c = 71;
      {6'd41, 6'd59} : c = 72;
      {6'd41, 6'd60} : c = 73;
      {6'd41, 6'd61} : c = 73;
      {6'd41, 6'd62} : c = 74;
      {6'd41, 6'd63} : c = 75;
      {6'd42, 6'd42} : c = 59;
      {6'd42, 6'd43} : c = 60;
      {6'd42, 6'd44} : c = 61;
      {6'd42, 6'd45} : c = 62;
      {6'd42, 6'd46} : c = 62;
      {6'd42, 6'd47} : c = 63;
      {6'd42, 6'd48} : c = 64;
      {6'd42, 6'd49} : c = 65;
      {6'd42, 6'd50} : c = 65;
      {6'd42, 6'd51} : c = 66;
      {6'd42, 6'd52} : c = 67;
      {6'd42, 6'd53} : c = 68;
      {6'd42, 6'd54} : c = 68;
      {6'd42, 6'd55} : c = 69;
      {6'd42, 6'd56} : c = 70;
      {6'd42, 6'd57} : c = 71;
      {6'd42, 6'd58} : c = 72;
      {6'd42, 6'd59} : c = 72;
      {6'd42, 6'd60} : c = 73;
      {6'd42, 6'd61} : c = 74;
      {6'd42, 6'd62} : c = 75;
      {6'd42, 6'd63} : c = 76;
      {6'd43, 6'd43} : c = 61;
      {6'd43, 6'd44} : c = 62;
      {6'd43, 6'd45} : c = 62;
      {6'd43, 6'd46} : c = 63;
      {6'd43, 6'd47} : c = 64;
      {6'd43, 6'd48} : c = 64;
      {6'd43, 6'd49} : c = 65;
      {6'd43, 6'd50} : c = 66;
      {6'd43, 6'd51} : c = 67;
      {6'd43, 6'd52} : c = 67;
      {6'd43, 6'd53} : c = 68;
      {6'd43, 6'd54} : c = 69;
      {6'd43, 6'd55} : c = 70;
      {6'd43, 6'd56} : c = 71;
      {6'd43, 6'd57} : c = 71;
      {6'd43, 6'd58} : c = 72;
      {6'd43, 6'd59} : c = 73;
      {6'd43, 6'd60} : c = 74;
      {6'd43, 6'd61} : c = 75;
      {6'd43, 6'd62} : c = 75;
      {6'd43, 6'd63} : c = 76;
      {6'd44, 6'd44} : c = 62;
      {6'd44, 6'd45} : c = 63;
      {6'd44, 6'd46} : c = 64;
      {6'd44, 6'd47} : c = 64;
      {6'd44, 6'd48} : c = 65;
      {6'd44, 6'd49} : c = 66;
      {6'd44, 6'd50} : c = 67;
      {6'd44, 6'd51} : c = 67;
      {6'd44, 6'd52} : c = 68;
      {6'd44, 6'd53} : c = 69;
      {6'd44, 6'd54} : c = 70;
      {6'd44, 6'd55} : c = 70;
      {6'd44, 6'd56} : c = 71;
      {6'd44, 6'd57} : c = 72;
      {6'd44, 6'd58} : c = 73;
      {6'd44, 6'd59} : c = 74;
      {6'd44, 6'd60} : c = 74;
      {6'd44, 6'd61} : c = 75;
      {6'd44, 6'd62} : c = 76;
      {6'd44, 6'd63} : c = 77;
      {6'd45, 6'd45} : c = 64;
      {6'd45, 6'd46} : c = 64;
      {6'd45, 6'd47} : c = 65;
      {6'd45, 6'd48} : c = 66;
      {6'd45, 6'd49} : c = 67;
      {6'd45, 6'd50} : c = 67;
      {6'd45, 6'd51} : c = 68;
      {6'd45, 6'd52} : c = 69;
      {6'd45, 6'd53} : c = 70;
      {6'd45, 6'd54} : c = 70;
      {6'd45, 6'd55} : c = 71;
      {6'd45, 6'd56} : c = 72;
      {6'd45, 6'd57} : c = 73;
      {6'd45, 6'd58} : c = 73;
      {6'd45, 6'd59} : c = 74;
      {6'd45, 6'd60} : c = 75;
      {6'd45, 6'd61} : c = 76;
      {6'd45, 6'd62} : c = 77;
      {6'd45, 6'd63} : c = 77;
      {6'd46, 6'd46} : c = 65;
      {6'd46, 6'd47} : c = 66;
      {6'd46, 6'd48} : c = 66;
      {6'd46, 6'd49} : c = 67;
      {6'd46, 6'd50} : c = 68;
      {6'd46, 6'd51} : c = 69;
      {6'd46, 6'd52} : c = 69;
      {6'd46, 6'd53} : c = 70;
      {6'd46, 6'd54} : c = 71;
      {6'd46, 6'd55} : c = 72;
      {6'd46, 6'd56} : c = 72;
      {6'd46, 6'd57} : c = 73;
      {6'd46, 6'd58} : c = 74;
      {6'd46, 6'd59} : c = 75;
      {6'd46, 6'd60} : c = 76;
      {6'd46, 6'd61} : c = 76;
      {6'd46, 6'd62} : c = 77;
      {6'd46, 6'd63} : c = 78;
      {6'd47, 6'd47} : c = 66;
      {6'd47, 6'd48} : c = 67;
      {6'd47, 6'd49} : c = 68;
      {6'd47, 6'd50} : c = 69;
      {6'd47, 6'd51} : c = 69;
      {6'd47, 6'd52} : c = 70;
      {6'd47, 6'd53} : c = 71;
      {6'd47, 6'd54} : c = 72;
      {6'd47, 6'd55} : c = 72;
      {6'd47, 6'd56} : c = 73;
      {6'd47, 6'd57} : c = 74;
      {6'd47, 6'd58} : c = 75;
      {6'd47, 6'd59} : c = 75;
      {6'd47, 6'd60} : c = 76;
      {6'd47, 6'd61} : c = 77;
      {6'd47, 6'd62} : c = 78;
      {6'd47, 6'd63} : c = 79;
      {6'd48, 6'd48} : c = 68;
      {6'd48, 6'd49} : c = 69;
      {6'd48, 6'd50} : c = 69;
      {6'd48, 6'd51} : c = 70;
      {6'd48, 6'd52} : c = 71;
      {6'd48, 6'd53} : c = 72;
      {6'd48, 6'd54} : c = 72;
      {6'd48, 6'd55} : c = 73;
      {6'd48, 6'd56} : c = 74;
      {6'd48, 6'd57} : c = 75;
      {6'd48, 6'd58} : c = 75;
      {6'd48, 6'd59} : c = 76;
      {6'd48, 6'd60} : c = 77;
      {6'd48, 6'd61} : c = 78;
      {6'd48, 6'd62} : c = 78;
      {6'd48, 6'd63} : c = 79;
      {6'd49, 6'd49} : c = 69;
      {6'd49, 6'd50} : c = 70;
      {6'd49, 6'd51} : c = 71;
      {6'd49, 6'd52} : c = 71;
      {6'd49, 6'd53} : c = 72;
      {6'd49, 6'd54} : c = 73;
      {6'd49, 6'd55} : c = 74;
      {6'd49, 6'd56} : c = 74;
      {6'd49, 6'd57} : c = 75;
      {6'd49, 6'd58} : c = 76;
      {6'd49, 6'd59} : c = 77;
      {6'd49, 6'd60} : c = 77;
      {6'd49, 6'd61} : c = 78;
      {6'd49, 6'd62} : c = 79;
      {6'd49, 6'd63} : c = 80;
      {6'd50, 6'd50} : c = 71;
      {6'd50, 6'd51} : c = 71;
      {6'd50, 6'd52} : c = 72;
      {6'd50, 6'd53} : c = 73;
      {6'd50, 6'd54} : c = 74;
      {6'd50, 6'd55} : c = 74;
      {6'd50, 6'd56} : c = 75;
      {6'd50, 6'd57} : c = 76;
      {6'd50, 6'd58} : c = 77;
      {6'd50, 6'd59} : c = 77;
      {6'd50, 6'd60} : c = 78;
      {6'd50, 6'd61} : c = 79;
      {6'd50, 6'd62} : c = 80;
      {6'd50, 6'd63} : c = 80;
      {6'd51, 6'd51} : c = 72;
      {6'd51, 6'd52} : c = 73;
      {6'd51, 6'd53} : c = 74;
      {6'd51, 6'd54} : c = 74;
      {6'd51, 6'd55} : c = 75;
      {6'd51, 6'd56} : c = 76;
      {6'd51, 6'd57} : c = 76;
      {6'd51, 6'd58} : c = 77;
      {6'd51, 6'd59} : c = 78;
      {6'd51, 6'd60} : c = 79;
      {6'd51, 6'd61} : c = 80;
      {6'd51, 6'd62} : c = 80;
      {6'd51, 6'd63} : c = 81;
      {6'd52, 6'd52} : c = 74;
      {6'd52, 6'd53} : c = 74;
      {6'd52, 6'd54} : c = 75;
      {6'd52, 6'd55} : c = 76;
      {6'd52, 6'd56} : c = 76;
      {6'd52, 6'd57} : c = 77;
      {6'd52, 6'd58} : c = 78;
      {6'd52, 6'd59} : c = 79;
      {6'd52, 6'd60} : c = 79;
      {6'd52, 6'd61} : c = 80;
      {6'd52, 6'd62} : c = 81;
      {6'd52, 6'd63} : c = 82;
      {6'd53, 6'd53} : c = 75;
      {6'd53, 6'd54} : c = 76;
      {6'd53, 6'd55} : c = 76;
      {6'd53, 6'd56} : c = 77;
      {6'd53, 6'd57} : c = 78;
      {6'd53, 6'd58} : c = 79;
      {6'd53, 6'd59} : c = 79;
      {6'd53, 6'd60} : c = 80;
      {6'd53, 6'd61} : c = 81;
      {6'd53, 6'd62} : c = 82;
      {6'd53, 6'd63} : c = 82;
      {6'd54, 6'd54} : c = 76;
      {6'd54, 6'd55} : c = 77;
      {6'd54, 6'd56} : c = 78;
      {6'd54, 6'd57} : c = 79;
      {6'd54, 6'd58} : c = 79;
      {6'd54, 6'd59} : c = 80;
      {6'd54, 6'd60} : c = 81;
      {6'd54, 6'd61} : c = 81;
      {6'd54, 6'd62} : c = 82;
      {6'd54, 6'd63} : c = 83;
      {6'd55, 6'd55} : c = 78;
      {6'd55, 6'd56} : c = 78;
      {6'd55, 6'd57} : c = 79;
      {6'd55, 6'd58} : c = 80;
      {6'd55, 6'd59} : c = 81;
      {6'd55, 6'd60} : c = 81;
      {6'd55, 6'd61} : c = 82;
      {6'd55, 6'd62} : c = 83;
      {6'd55, 6'd63} : c = 84;
      {6'd56, 6'd56} : c = 79;
      {6'd56, 6'd57} : c = 80;
      {6'd56, 6'd58} : c = 81;
      {6'd56, 6'd59} : c = 81;
      {6'd56, 6'd60} : c = 82;
      {6'd56, 6'd61} : c = 83;
      {6'd56, 6'd62} : c = 84;
      {6'd56, 6'd63} : c = 84;
      {6'd57, 6'd57} : c = 81;
      {6'd57, 6'd58} : c = 81;
      {6'd57, 6'd59} : c = 82;
      {6'd57, 6'd60} : c = 83;
      {6'd57, 6'd61} : c = 83;
      {6'd57, 6'd62} : c = 84;
      {6'd57, 6'd63} : c = 85;
      {6'd58, 6'd58} : c = 82;
      {6'd58, 6'd59} : c = 83;
      {6'd58, 6'd60} : c = 83;
      {6'd58, 6'd61} : c = 84;
      {6'd58, 6'd62} : c = 85;
      {6'd58, 6'd63} : c = 86;
      {6'd59, 6'd59} : c = 83;
      {6'd59, 6'd60} : c = 84;
      {6'd59, 6'd61} : c = 85;
      {6'd59, 6'd62} : c = 86;
      {6'd59, 6'd63} : c = 86;
      {6'd60, 6'd60} : c = 85;
      {6'd60, 6'd61} : c = 86;
      {6'd60, 6'd62} : c = 86;
      {6'd60, 6'd63} : c = 87;
      {6'd61, 6'd61} : c = 86;
      {6'd61, 6'd62} : c = 87;
      {6'd61, 6'd63} : c = 88;
      {6'd62, 6'd62} : c = 88;
      {6'd62, 6'd63} : c = 88;
      {6'd63, 6'd63} : c = 89;
      default: c = 7'b1111111;
    endcase
  end
endmodule
