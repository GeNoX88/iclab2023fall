//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
o7ST8oPOwgIjRPvfBbB4nyMb8LWuxdYyVZ3y62ZqrtygSad+sLVC5Pu4y/zkZCtl
gliXaWrxsWqh+cDIZqjAvVlePV8ZLrg8hXXZsm5ZZBGaZUwC2X2KD+SrZR54hXD8
ffvqMy9Kb+3/29I3S9BODpmkaZMhSKkt0hZkXSrFOmU4jgnsa986tz//tGkYHcmH
mXh1s8g/twV4OdWOkHq5i9SYAHmxdMFI2hfk1PkKJJsTQreQe491rKiondVmGmcZ
eoTQOGNLEElDcHS29fs0k6shPJ2p8WTn4wiVnBub4CPbq5/ZGfhBAKLa6F3PX/lA
atoA1huGzPOIeeObI0bNsw==
//pragma protect end_key_block
//pragma protect digest_block
9O/wCpYELIkC8dMgvWRy17tksl0=
//pragma protect end_digest_block
//pragma protect data_block
8Xr6UNszQfTtS8aoMyXzujt//KoMbz9QzdJJoep41jiZSKIIYalGWn8h2xNohH15
M7e6KnwteSigP0lOSZ8toTRiYnOSgsROWzfnLuGPV8eL+tBjho5Dw6NBUQTKicz7
B8LnznQ8YqiyQ61nwXMsd/JAHqvpEFLW65wGkjnI5+cmo9aaUln6rljo56SBvkaL
yYt/595YkBcI7NHzwAkX4ZGkqJd8B+MgHOz7LeozerqdBlUFDBWHnLwNTav+lwgA
To/Ci+fAFEbyVtc8LfCDfml1MAzvT3/e2jg0hdHuJX7Rbw9uofT85LCf73KA/kL/
ytz2np2neDpPUxlxEdPctt3tqgk9TLp4stpj/viAQ2S7f2/R0HvlT83pFps1E9f3
4wXNusFZ5fVkQtFpEnsCLgMKS19G/PAHvjOliXzVqmwqCzU1qa+a7CnPUn3+yuba
WiWV1wP3P38FvM2V1ibutx9Uoo8Rq/676vMl7Jv5qf3XOBeqJbI6d3voUW2ZmwNJ
aTniEroyUo9rwoM4idpjoP70GDACkWvCsNnQJv1jlTYbVmRfH3AfP3226sqMbg+M
uDDat1FPzrG3tH9swVp7PmTYciW6kIqlAs2XDCgxzPM3yH0Pe/ZufWyh6fgSK+cR
GAChoNFs65Zti9irpF+jGLutcaTJyOoU4FY41Cf2gMz3Zpynq/8yibTSXNO9hSEM
GIm+LdMUK7J+y7WE8zcuiEfjkIPGF1ASrfGTYKNP3YF4U/ToGs9CKPB3VKMt1lIw
fUj6TppQ04WXi1pCUa5AdLAUA0sJVfrW2PqcGueuhjiqQizyaqZnZJH4hD/WFQOQ
TZGjdmEFHJrVuw2GMyOSSHhEQ2rYDDIT47JZwDxP+WtsaYv40wpyLAZdm7cXzX61
nvlQcOrqLkRjn0iNaQaPNWha0GW7zSAVYC7CGtHqjs236fDmFQRLvimLTCQSxYJL
7G9lLimJTaCyamy1/LO+YuIy+aUTcUA9Q/1H66M3Fb/B4mW3HG8lf6CkLKjgR/NY
wb7T5vdW4IiJpWeFXJOoaWfMr98XCiH4aQBCz3vyQbv+gPRuLGhkozTJ0Rql6ppt
wTFAWQT3DWF6LTcu/aokSUWIYDds9eCCs+IyT4OJGBCiu+r/2Gnc3fe1I9RydtPG
PtVSGGV0uRSq5w8VHwltIkl2SRQ6kBCRO4F8UNVKT7cpw+gDDrymul3fJBAzEjty
pBMpcrMUc45Ykkz6bVCce1wxIM0MuJrJTnNcZ0OZCwTCCUs2ndKaTsfuVUXYqKF9
NzPTvLKsvPdKnw7dfyMzpC/3+bV51wHigzi6PImzcXO0FpVf/mTLLxYzT/b0QkIa
8pBgFLf7EW78XsTJzwCi8SSLSCQxuarpI8fynCosodrhKc3ldOlNhpgiuy0wzSUV
ziZrTJUL4cpkI2dbGOj+zVdfbr5xquYCop++h1hfn/SQtzdfOJfctxo5QtMpvkSV
FSU2kZicjOUJ5eby7TR1DdNtlEhd0d6prxDsFOrDft6UKfqKFyEY8Eut7W9YZxqu
4APxa0B059cf89LF7Csg5iwGaBfr24ShKDQDq4OllbmN7XhL0fHrffbfKgtFpJHQ
PWN5u93ylWgdiKyJeb9jiwbE0jYoE6JlyrvHHrs1q87L7llbXgVJcn8PzO5+y+Nm
ZJqoxjt1KigGxn+AvBoznMZ1Ddb80CJ9AiQl2V6cGCllglaY9Ck5ABCPzEIR6PZX
YbJz/8rmHnG1sn+oeLUeLp5E5jJxUaovmsOPcEqjZMnIeC5nfGSd8rQJNohQPvi2
r3ZAtv/ovXZ6G47qu+rvqfy4g0Yo81CRgU1AiimEFv3o9f7h+jYc2pX8KbUU0+Sb
ASA88dJq//SNO8peu3I/Hqm296NHAyHWqCwFlZHwKkLivkWhA/wDWlldLAOOKzBe
/731vfYck9s9bLCnVM7vEv96fHkZEESc1v7p07Q0AWP813w1byPXfsMPWn9HQ2ps
lL6ZRRQ1QN7XTXksFNpcDyLK1dzu6vQyw+cEwH0aNitRyoUVGLWZ1Svaw5sD2pxH
jzxXeScZrWg7TJ610Tu4ETdo7abaq3Flpdx+DutBSBCk2tCezUeB8nFAGuSG6B6/
yFrqnm9GDi4glCWBzewBQaK0J2+H1tVnx2SiGGWU+f9DiDEUSNVArf43HwQuTUAk
DK+9vgMAf/W91fu5RjSt/K5DVJqVofPWiwdhyie1RPearYT3V7LW7puWJNweWfyZ
nkuagkld7MKVVi4ZqnWjbYq4XTTB/lL0VDk4WXsg2tl789jVAqKOVk/q6EocYMua
uQUX0rapIGXSZsTwZkwFsJLlTp1ZU34JXgFN5YWf6ULYVF0Z1pc7CDpyd3vp5S9S
8CMHz26HtM1VPy2f93PppRtIWIeXolG+T042+i8PMIV3Uhn5QSewPcbdm1RzuHCF
Es0+qNzFPUhggch9AhUvSsV1zGrRsfwbbRXDheeRuge/66DnJBgM495H2JXyCmUv
B4Kdv2QIDj5Ia5wgUWs7jXIBiJXrm2x/tPR3g9Lsn9nzq6UHiHR0Oq6YS//0lMnt
pkf+PnVGkfoHXhnd0YDU5eb1Ru14pvFTE1hUwgdQ4J7cvXcNVnmEzHEqT3s8VplG
d7xYyBoMnO2Nn2Wbe+ZaZugbgXhSfBbgwMOlzdadaVjcAxUlU6SxunTE9Jk4JcTW
qWA6LcaG2QtqLErA9X9ifl3TWIRfsrX/dZZaYimT8PmnWudivyzqfM929gj9HPjJ
aAKyELrXew8HwSwD4TLzbSvkh3z5rYJ87AqcMLSYnmvfbzati6JffjqxNvxGjncZ
Y2OqYnbwiaH50I8+8X3DUgIWndUx4xg1Q/XTISojstN5wSyFhvv906h2rJCLKNwB
RSiejmEPkKPRv7Vo5MxlIAarir3N1kQ+UlIkfi13YbyWgnrmkQjDpcrQEud4QbEK
uK3+Uo+gIIKyEAwb/2jT2KnTK8ej2vD2N3cyMrWQaYK7oh2kdBdhiivJgfth977E
5IzAOcR3U5CQ62X07UcxftzJiNGaXXM2V8MPhlKHMTyE+kpUq3z5iVizmTc+ADT/
ZveKOYxL1Ry0C6IgQV8Ee5QWA5UQiogxgP+S41yHtrrbKmL6dDKS+4rIPaXBJv97
luBt076nk38zpJNzNv4r15Y3bRqrhQcDR38RHj4zD61RsO/3lwyjNjPdUS3/RkjF
k/Q15+HX9ozc91vNGQZzEOwRQidJT1908po0MygxlZLWygI6txDg5bOjbwkoux/x
qS/OI9ZbEo5Ki8JYmSc4ELW3ScfCB27K3ar0EINXxD5wUQXcUslx0thm9Ci4gszQ
NiDcZUDL3nNpv7VmwvbjiBQ1ISgvdBvTF52DGxtPfyF8LuNZlBf25J1LD+k1bXLT
NOmGVSzHx0rf2keWloW59Ca46UxrWnhxSAuCKsxIgQKRJftgeqJlvHEJ49fUU08e
kVEl3EVC0OZ3ADsphXQzoC1BInN53QL15EUxuJDB2fhYJtX6ZcCHRQU/oJJt8CAC
oy0ABnOCftUYwQq7kkKId0qNGE7/jLBY9X0Sj4GWrRj/9BKhlo2mYbg1v5XkkjQk
eMyx4lozI6J1UtnLQuWLukH9p6SMV/veKX/Q0lAqjg3yOj74JZUKRf6AGsgwzQKT
7hjCmN5adqZBXtbwzH3uyZmIZhO2j0/uRtmwk6oiLsHENdZ3eyahkd/XyFWF7xcR
kDle8LOP4+JfRRVqqFnifVfsDFfizQSZGeUXqevAfVgNN+quiem+RwHCnYbgxcS9
ZyWi+t/mKy3RSScZRu2csdep3v3TXNprxPKBu9DbktMo6dPhAtf+UaE6AC/ys28I
hUveAd/oJJ3h0U8TWqdA3xXGjx5/kDXjurthSKfSrDEGXkQS8ky9+rtcYExiZM+2
dobAJ2KuSyV1okSexNXZXTSylq2ZmVJxsaQBHwWEBFkz6EI97BGWk2fAiE/Ss/TU
AS0TNoT8AGTbwIhTcat+KSnv7UGYQAsG+d75ztCXOofnIW3mVm4xa1/S9b34eQCF
/OJjhenPpH35Zt82YJhnPShMRyBZWTJdQ2kTZ4yXng/T80G9ACeNEs8B/HWkaVuh
i72ZlE9v6qyMRcvgdxMCmwVX55H7npSCTbUb3kf6xzU03cuX2Hdism+ltsAcL6Sq
3m3hWTp6CfJd/RkH7jvewTqh0wVDR7rbclbz38k0jHa1f0J3OdtbnT+mYiXQjbbQ
a76RSUhTjF+7ULUqEQM9UNhLn+bG/Zu8ed7Lkl5f8oM7YijGFanEROq8hvAnoDfy
SIxCxB9DqS/BmpfdYpNUSsz94ppGJW/XqwebJ22qd+Xh5ejWp18XOj9dAV+miIpI
nvjL7QgS9MEcs6J7/DsgFc4Pp+yAzcO+vMHEwEirmyYuRGi+kHVxeCEG/Tus7tNE
vAOLHJ5EFNde4lTMGYsya40I6vBYnuXcAPtmfLDP+7GFlm1qnzJ+lHbUZKn3T5HH
HsuCFOXe5oWBnrAJFs6yahVC7P0dDpcs516gawafGqUsfgYo/6TCNDnV2+E+Myw+
JbOG5q/PL8BuW25SGmkmxioCHXmRmX56jE/MwEf554jHcffH3NSJrBjsOdpgigmJ
EZf5PgjKJ8skq7F5dWHsAmut1ltbHYV6k2nZnNClAE3T3KGn2DpKZWlkJ0HVeQq1
1ZQjfThxeppGgj1OZxXjOhMegr8ExsPpF6hTPsE/Z5Rspqp6pqpoIhE4v7qwypKq
K84m3oTpdawklVKxra9OTmGIUL8SFIwh2Ur9CQhJwDcZb1R5RlU+1XSORJthQ1Vx
XDh5XDVOuzqBlUO9PlFRo5IVe8jdC/eb1YGidM2kmwF4yjsANx4H7G7OwYfdf3Tm
F2cRQzOdbnRzmZ5KEusYzEBkGeoRD+YivWpGZopU0FSdl7a68j3qj9VhONhVsfun
a0hrbNvpDBLDkePQCXx5TOtdeIF1kJVgzAUcpxzsGjo5+bTXapvPFAamKBvaJOFH
WrPydjTRMquWGp1hppZ7FEXPsTDd1ov/fM6aHILGqgPTlDHf+E2dy7LBV8ZtOgGf
ypVMxM3yl+t8TCgJCvsrNZR3yZVLFNN80N+V04IHTtlYac/+Teu2QD7+EAOa053C
qK7ehQnbal2eF2484Uf+g5hv6XmHJP/8yBAC9r5N93Kmrca26+CH/OKFVdzl2sMg
AKyv+rhEZNOsd41REYZJYzbndjaUSSBdcoGQwXtL0xUXOkPg2XBp7nzJpx070my0
4M8Nkm8ItV52IbNADW4riSONvJfyMb78e0luVPKCTjjIbpRtxvLCI2pKlWaczW6A
+iaKYH6h7VWE1HkG2MbU3tVRRxq/G8rfgfZDydqG0AcBRQzBYE2qaz0DHsJgh9G8
TViKnCxW6BQD/iIhTbrusCeK+AIeAEJ++q7QgZTnYGtfD6AHX6nHkujO41OVesa1
MW7kh0jvqm2iHwIIsB9OCQR058vmNMr9hISS5/ytFzsWrcjLzaexVMy5YbYQIW0F
jYWsDTg1hW6dI/v+AM9xGI0+bE+Sf/K+G25cblfyX9cOTDc8s0qs1rkyFILpybUW
HOTOZN0UBFWhCpyUEP4rNEWd0jYGNmVye69Bfdb6BnKrrg1tbYhj1tSLj40jFbtC
iwAjkwuNu4vJWK3Y7AmDukKRY/QPeO0Gqb30Pa8nEt/iZecFLEvvHYXQEKLTySJN
qEd5+7msS6cR+Oukp4S7OGVwws0ILdELk2yiEnX7apFmyxAnmVi6hBbsPHg2qUmp
t27xMDLxxz+8Omn1hsXIintVhlAqNs4CEHloxfKCNYXL9xpGcYaMi42l0LEW6/nk
GjmtLwOiKJ4fLOIQdGPyGQUOvqZtmRcCLCqVNC02xf5+SAx3S64KO5xc47eueIG6
ZsKcbPtLaw9UuJWVx7m1O4b/AhxDI+Y8zHxQCZcDOdHmj11yn6CEPqQwuf8rpm1z
rH8JMeR/i6OnjPg9qCUoFxOYq1hR9eKjoFrSIlmd8DHNbaHETU4ym/x4MgrelusN
sy1QeWU3lNcdmBeT8CPov7p/qks3lUQkzxzD9pwnSToA88rFHtJYAu80s4gOCURq
0t+Do8xpyKkxLkktce1yzxogNlQ9Rq2q1VRkDqC9FmZ/k0jAB7YGfEN9nGLwIoLo
8y6PZgfBd3llE2eJk09pQxkbwZgjL7waWWHQf6UQyCTKsDtBc+GeNIzV5OKKWfcM
Ja8MadBPCYLGvuvEbJ+bogmledhKertzgSZxWKWK/RA1rmV51Bd/uQhSMjJ8iZlv
CIQq6VH6NUXBoq2G+rIlPaMnoZ6cuIQStfOqS/PtIWznJRZOm0ynomqwIODnRsH6
0gMqT14qT/dfbvBySrB5O5Uj5Pu2tPHND91p70iUToMOdFCtoQx2LiLTa/quGRVe
lsdvvFf0T3UxFPsr/7Wd9Mvr/fnIfsxfLPVH4jUTeZJ2qCTSbLD2GGlbpV/9kgs5
IFMfIOyg+/yhPhBXSjQhdixt34mr3WGKFLc6iX03W/eeenieB8xuauonxxMNJaY5
9paJaCx72muJ093QeuTaKaZRqMe5XfKcVp4cHEm07vrwe81NPwnXOfxo0+dc9xlh
mgS1uMKCGWFwHW4jd2+YBw55CE72fQbGWJPl6eOWyY12UFqMqBmAdqlyfFXRAhJP
xAYyWxj2GrJUq0+2YwZ1TplrcEPveUCK7LF5p1tdazvFNoJMy/S2bnlHGFt0mCQI
UwcMTCoTTXuUl4+EDIdX8sYtnVhkFE/OAT/yPl1/4zWPF/kgZDokyyANgEsC/nrs
T+Pct57V7wWvix2yxvZqq/+EzcOnm2SkxhP/e0GfidGSkNUf+SHQFtxAuu6vjlI/
OJXfOPb7283lmBC0Oa0fvk66PRfp2oyQwagW5rcZ9L25or5k+eK7zfJEogx4Oucl
QPvl6DRTaMxk4yEogB7IKUET2IDfcDfIMj9TruILG+4HUiQtwgiqmxH4sUvXOueL
c/CBvZA+LQTKei9WNS1KJFLw4vzNxhphZ7QwJm7VWjnCSrRgURwv0SEKGVrYwAck
KF4V8QYeYSHkd92d4Zkvly4gMKlzgKVcDIcLwcehPsQoKg54FU2Chqy8GW++UVXT
ZTrItKhdQuS3nkuPfcHqYEVv01R7Ag4EBHFTOwWJo03MzXzFq0yJkzZn/8+o3uwt
To/gNbPFaufyNztfigogOak84cESxLST4j9oPWMkEw+4RSjm54ASkcC9XKvIH6YL
MsRnDFhT/wfPvR9/599oLN2B4ka+J2zdnJ2mW1kGc1moVu+iXj6E/5PkzPYejGmF
J1pNKjFQ6DR+CCnCqnEz9TuT+n9jomzvUlN6vOJjCwMuItfYwK/tuGj61BoH2fMf
DiD4/OUkRzP9wMfJqoTi5inJSXbRQRUkUOyj59sSbqrp+I2q2ET9xcUFi3sGCaNH
NAgPrAnsNry+1A1Y/aFbneKWekele7YzPyw3AY7aXJ4F7tDM+D4n6fDzfY1zvOmh
z2RirO73mk0g62rt0UAF4v/F6VuWg3VXH1tySLs9a8xR9oXqS+mzAjfjHB0eDgps
hSrfcvzbk0huZohTqDzEWRmAAS9blGA7D5FAhyfqwcovZYXb1zTLjf7ukHKZQjx/
EviO68pO/K3se6lLv4whVnwlA/FLT5a6hzOjZh0D/ak8C3NTYGtOB0BerKvtF1oF
ttkrEObAUc3VRoiQ4l2dT+/PeS+k3wxt6EdxhBiLmw7qbyGYs86+ONxxKFgukYqr
yxaIJrcpHu1M2cKHa0fp3jfbVNW0HrYjBf+FPSjM62wtdB1hJIbjn6SXKFVXlYZ8
IXRHs1C46l3jo2U1BEd5eYiQU6Ws/xxAuB0w7C/yU8ruc2IZTumN7TobgYJJhQJ7
scaFeoMwf9sSgnb3H134fb5KkQ03AOFF9f0fGvi/7zRrbxC17UzW9mQRjGXz6SSN
Ew7rozSRhfLy2rVnxjIWFqtwsIgHW7X0FB6aygv9CS9TB6d3Pqqv541Zh19h6dJD
xvnZRvI9ZfZ1AGxhEEOTGucubHF2V4fWxp8EUxkcbhy0+mCVN62OM/BPA2BvAQFJ
qF+l5OSxSFEIdEk27ODxlS7zpteOFz+E0vlkcHAw3UO24CwhAneAVKH9gKkOg/h2
rDqzY4bcF/rFqK1bTpRc8B+shr67ojjcgoGvd11a9uHa+bsK5FRxKRcd0Imoa5ZA
67JjwuHz/pgKinaCsnn8xrsfNSAzVgMJ0bc59VpmjjDHY0SSXzFcNrE7TLl3sDVE
8nQVuXd8TaUW7S2IAC5XUdtWc0TBJk7Y9N85zMkB/ux/vqzP9iLyu9upUPnyrn6b
ggbdaVmIWBJkwQjOcLhny5bUfPsijsmS5E0lToZH254Fcqr5zyM3vKMA5gSPn2aM
R5auiek60lK9dXm1s0Ml5qQMa47DFQztUub0MKq2SFrFwx9IxUmwO/E/r1SXRRcp
HHJUVWaP+UBEdeNeYkD18gy91vyPYcDpSUJNJaQMQJXZlWaqkum3/jnC5JG0ETdd
PAVvlumWU3suOzqwYTZiVEiobbmM+NR0Xh92rQLEzt4T7Ocp/6itnirmbbOpiJgp
XwYSqFQQ5LgM/NCtqFCb0lI2FCMUH69/YKPe5coy5a0kjbL3BTa/m1oOWR4x92Wm
UesL8il9YwInuTGcLsheCyoleEDsV4Ghl4ERAposk+PMs/9KevrmsYNZ79tPTXAR
caZu6pHFhoF1eO/riG7JpmMvXp+TCgZCo3smd+XP+8wI2BiqNAEEEEuLFgYYlTFP
9Zcisr9oSMf8F+C47pF+TqYcjaX7TYwDVtNqN5i7DxaGghtNvr66ZsIPBO9ihMIB
GvVOLzgh2IITt4IjAjVhxgRF+vhxU3ECoqzcK7It7ViLQmoID7/glBXPczIuZ1Vo
jnweoGtPIo3+cm6LcFWRpWu2j7jGY9R4w+Oofkg0OAyYn21Mv0VwXeLvOpaV9wUh
1xrFq4zfXC7EfwYwlCdjsejm1LPlYlDdPsKn8IJBwbafCBXLFeBiyMAP9amdu1LM
eHQefRLg4sBvn9yoLwVOSHe53vI6IWdbxksii+CAREqw5kruRTZ2EW9b5nChujTN
2+o83UujGOMUsBC3gMPRJIczVcX7RDu9yOtivggRoWrSS1iG7+CzBMCq1JGcEWWb
4UnXH1HIysTio01/hP4zqYXEw5boC9nOB5ZMtd8PUeqNODUsDX1JeuZ1GYCNdZTC
u4+SoPxz60dJU3IE5SeztKNDJJTCH4TO0qctWZC/zMe72hw9B3xWfcHejaqgwNDI
B7RoXcOFAOA2G/LokI8QEnn2YekwQxbHwMMKljl78bU9lsaWicw7JBgG3zTsrsWF
+uVlwbQjk6WQy/N0JnKFKnXcpQnmr8N5e7VjQcY+ZLULS2rQcQYcZozMsNj3D8gg
/4p9x5tMIFVuIlI78bwb1ASS5VkrpbRrzSvnkxId3DfvZMOJFTbc5XtVruJ3dYo+
WmdtKV1+v/FW1MiSrmkBRtP6vaFhAnYr6hh/spmsShPg5Fo+78ZZMBIi2ktwcikf
eL+71kVMZj6liGjmVIBnDn8nSwdhzAapo15yGsXKiVZPBnZqOFTyxjMsyhpzXOCy
RTIdEW9DgIOJdHmLwCT1MO84PUwdW/UQMHBYHzTO8aWYuqsI6hTWxeY2fkWyCOI+
r8fOWQUkLsAj4/47ZwSwNO24dAv1YOz3nDdwrdMPWMI3+IgOlTxxwzFCWgwl3xs9
1kLHKVm4HinZTtrBp0nZVDTE9dX2XUmyqQpbiVrgaHoSs1EvDrcZc9IhTuuKwseu
NzjgRxHf0cHa8KNJrEE8prxYsheeragc1VCk3b03jf9Es0YatjTPWJ4kBX97/9wv
G6piBRNUKSQM39x6VLSWTcg0c205rufe2XjEs/nkz+VCPKPDJ8lbR1RxbGcl2z3A
mKBJSVcQ/feyGYxIO/4WL2JTog1LO1WN2yF8imrf/BmOKPDbQCUKaTXVJ6GDinNj
ggVREktLgm4UPQ6W/86znfLCH/XBdOVPHWYtVP5S05KFhW7ZwV1MnihUHsPzaZKB
IQWvKnALpgGOnSuoENyD3k5UHmczWyOCkihpKawS3XjvdK+1iSJxoTnurG2p/xAB
sfk1UiZDZ4hBEQBvNF3PSealQQIUoSMPbY0ybqGG8nofo+B0LOo8PcvKjZeIESXv
sSz6L4d99v4NnmnX92PCbTazXxCbQIGGyzOe8+oe1nMeOJOPeaeb3RiqMDbQdm3a
K+bdV8IkOTPTIWxjQ08AMMLLcnyq5rTvD7imK8GB85/w3xl24LviU6WsuqBIoWFk
iO1QSe0Q0m3su7YlarVOKVTS3QzyOcBRvZw3toFfurlmcOBqoOgUO+qX7pAxdZ/w
WzSvPXMEll8p3AgeuCdv7ZxcZ0ZfcewqJQqXz3EXYsuWVkPZ+ukXBvuoImqqQnUA
4ld2xOfSXMtHhLWPN88pgQ/4WWS/Sofj3duigJUCgUgB+WnqHbJwVDdzbxscbkLB
BsXc8OXcovfjrvrg+PmIbMuE+9pRqPnlJiqNs7CU9PBMymAJqlYDRm9MTVCE5OqK
CdvSV1wLU0ncc4rLgvzTSmDbmhZSNym3jYFxCdo92IA/HkKkj1gKPA3QMvSWJumI
PGybzvcLxkSaeZs09kkQL95KsQdzNP6rgwXenBorzx40+7r2JSMkwwFDkadaoSla
0jTuiuJpmOvJQtnq7Y0kyLbuAuL6kfmNVUIHHLDtKmXFykTzH8jkOt4MZQZpwLNr
oawCPnGpnsvfQmYdbHEaKYLpDngo/H3dixQqWfMfn/HczeXB0UgTg5xC6fFog1QS
Q7xzkS6rkiSMxJll6SItmSG2OtP1AiX5A51/vTmY+NsXdeacO/ko1IZFzSCc/Ceq
/5PP/s7Ayd3K0ngcL5MOhOKig/jKNtxpObocl+VsCq8bQaLj/XP37/WdcnNwPL6Y
uXGlXlN2/wRY6cqaa3pJ07qEDcjLnZ/DSRFM5aJ3FytaquM8NL08OlXc114/JLZl
Zjenjwwlp47eRdCAwIhyTDmBjZ1u+WUezzc9fNB9zs6RXXF2WPQuir5o1oTUE34K
9J+urcS3UAJ8NfBROSB6jsFKP8qlj26Yc8N1siho+RjPH3bOfR7RzZNb1qTHYzQU
8AFs8uGmwjzLURcOU9FCYah8fMCQwsUYliDWT2RI02Zq2OGtuKVWPvEUrnhjqnNo
cbDk/3c6VUahZoC/8L/0WoP/fjh/3Y5GBNlB47jymMB+8wHtfBdjs6T/pHotskyD
IqsRE3q5F0lxajnhJCo/jakT3i616Ic5CD5nV2zZnqE7mlUqMJqmqJVJ5feTKhqE
MIThnb5qUAh17vzjXC+bm41GYTLJim+5XzRECWv8amOG8YcmpxLXM7jEgVZYc/i0
LBW0lhXVUUVdtHdM329LrASiscpjxnM1vQrwJ/YUmCBXEECd4UQRR/74CRpXk4nd
+J5kmKZikJb5AQXHcvJvvvXNRy184c1RrqZHwHN5z5+DK2J20ZprWJRVWtuBpYLk
PeWze0z9BGnXrQQRR8/uV7CW0FFVkN4ETVK4MXZ1TT0sgA5l1yOQ1QJ7lPu421T3
logxoTGLa7ZlbwXLWknBEw==
//pragma protect end_data_block
//pragma protect digest_block
/APUl26SeKiwS8YVM/5w5vQsWC4=
//pragma protect end_digest_block
//pragma protect end_protected
